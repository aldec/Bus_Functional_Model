library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.numeric_std.all;
USE ieee.math_real.log2;
USE ieee.math_real.ceil;

entity AXI_QDR_CONTROLLER is
generic
(
G_AXI_ID_WIDTH		: integer	:= 8;
G_AXI_DATA_WIDTH	: integer	:= 64;
G_AXI_ADDR_WIDTH	: integer	:= 48
);
port
(
reset	: in std_logic;
clk_p   : in std_logic;
clk_n   : in std_logic;

ACLK 	: in  std_logic;
ARESETn	: in  std_logic;
AWID 	: in  std_logic_vector(G_AXI_ID_WIDTH-1 downto 0);
AWADDR 	: in  std_logic_vector(G_AXI_ADDR_WIDTH-1 downto 0);
AWLEN 	: in  std_logic_vector(7 downto 0);
AWSIZE 	: in  std_logic_vector(2 downto 0);
AWBURST : in  std_logic_vector(1 downto 0);
AWVALID : in  std_logic;
AWREADY : out std_logic;
WDATA 	: in  std_logic_vector(G_AXI_DATA_WIDTH-1 downto 0);
WSTRB   : in  std_logic_vector((G_AXI_DATA_WIDTH/8)-1 downto 0);
WLAST   : in  std_logic;
WVALID  : in  std_logic;
WREADY  : out std_logic;
BID     : out std_logic_vector(G_AXI_ID_WIDTH-1 downto 0);
BRESP   : out std_logic_vector(1 downto 0);
BVALID  : out std_logic;
BREADY  : in  std_logic;
ARID    : in  std_logic_vector(G_AXI_ID_WIDTH-1 downto 0);
ARADDR  : in  std_logic_vector(G_AXI_ADDR_WIDTH-1 downto 0);
ARLEN   : in  std_logic_vector(7 downto 0);
ARSIZE  : in  std_logic_vector(2 downto 0);
ARBURST : in  std_logic_vector(1 downto 0);
ARVALID : in  std_logic;
ARREADY : out std_logic;
RID     : out std_logic_vector(G_AXI_ID_WIDTH-1 downto 0);
RDATA   : out std_logic_vector(G_AXI_DATA_WIDTH-1 downto 0);
RRESP   : out std_logic_vector(1 downto 0);
RLAST   : out std_logic;
RVALID  : out std_logic;
RREADY  : in  std_logic;

init_calib_complete : out std_logic;

qdriip_d : out STD_LOGIC_VECTOR ( 17 downto 0 );
qdriip_k_p : out STD_LOGIC;
qdriip_k_n : out STD_LOGIC;
qdriip_bw0_n : out STD_LOGIC;
qdriip_bw1_n : out STD_LOGIC;
qdriip_r_n : out STD_LOGIC;
qdriip_w_n : out STD_LOGIC;
qdriip_doff_n : out STD_LOGIC;
qdriip_sa : out STD_LOGIC_VECTOR ( 20 downto 0 );
qdriip_q : in STD_LOGIC_VECTOR ( 17 downto 0 );
qdriip_cq_p : in STD_LOGIC;
qdriip_cq_n : in STD_LOGIC
);
end AXI_QDR_CONTROLLER;

architecture Behavioral of AXI_QDR_CONTROLLER is

`protect begin_protected
`protect version= 1
`protect author= "unknown"
`protect encrypt_agent= "hes_protect"
`protect encrypt_agent_info= "Aldec encryption tool"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
KWEx4d+7fQoKvRhJZNxzx5Edpb0RjIoiqP4EFp347MAhS/4+5rLeofroJLad0LopP0oUiAvG
Trb+8jqVNWK4Gx9UYJsX5raL+ijaJLK0fI0dH2g4fCSBPB4YYyDtHQ7ntpKlqByAHybrJ3FG
H7cLCQlA1rWI24KYxYNcc5ajkyvFmxBmfIqwziODGoUEpB1swn+TzFae/Jx/QKqda9iLvUBw
VRS0K8tbxBd9FSpezR1fF9oaD3FvhuuWpzNjefDvzbPnMe3DRk+22tIvZblgwh4svlqXxe5/
kMDm5B4XdXt+uCWnTrHlPtmT09Ya9O0co3o3Tm3pLvXfHV8RhUM8Lg==
`protect key_keyowner= "HES", key_keyname= "HES"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
FDlVyJ/XNsrYQr0wWeKNezbkR38SuV8qe49SI0WkmwWpnQcZ2zew8HZJhZQku446yp2QlOaX
85m97GfUlc02L17xhj069j32Zh2VoemULswZxkk3z3obEBEhtL5zUJ+qO/hog3clB8Xwy1Jg
VpVVyh7uX2TqaeIPCPrgwpNU+ghRSEoKfkcYORXApXwRwL2+9hG6ZiO7Lr/Spjz2WSs8A4mt
GaKKzm41/Je+ZHG+IpgLkIGGwwG2K6sxi77FPwNG6Ix4VvPvUG1opGTc6gdWzhHZjkSqwnx6
YYyIuQiMXcvS/C+eqrMrNRZrxbcxRGyA/lxiVk4VSsUw/xqed7HH/Q==
`protect key_keyowner= "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
RJpUcyw2hc4g+YTU52WRX68KgiVQLn8/Ah66bO8nhxx2sB/FJlTK5N3dir8KeDvACzN8sc0x
aF9aCvxnMwRdvKMVKpULfPl2bkbXAdBnRtRCuviDFQzn0lJvvhjCHhZGdTRAy49r2gUucsAM
xmpB+0+QcvafbP/GTIIjUskEiy57k4X5PXPR6z2jPRoZTBQnP2uDRhV6dGPctGL7NxPnRDfR
b6B+7YdH0rW2163Mzqyd+BNusKqkcWyKkMNP0RmU3WWMHqyWK4xKmP0tryPa72kgo6pDsBZa
an1klxuiG9KV9KYfvpAxcgXql1FmOanWLawaA+zl8IppW0BSgRy+5Q==
`protect key_keyowner= "Microsemi Corporation", key_keyname= "MSC-IP-KEY-RSA"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 960)
`protect key_block
BRoDRCNtbrALVpgst5+0Z/ix+wcFeMAVzvwx9FTlr4h8nB1unrzbhrmL7uqW5c8Cw/lKBull
j0mqYbEpQKyIKbikXCcoKFo3g6FbncurRFlAP70tyyX+X3SF7xSDy1oi+lztLHAVjKVLLoge
CKAIM2pEdJCpG/idGpTTPtQSJDfYHlCHobzjQ6WZqH0XWd+CSyGKy6tozigiG1IvF1vWc9z3
XRJXYVlqhUzdR+Nxfov2Dna+GJau8qujW8xkV8dM5HxA0rnwB4aXtQVPrDWBEBL2agV7dyC/
FnOCK1PzjL9YTcLXEbTLoDOXJn+Wo59o/k6l3pFk5901CEVuVmPcTJQ+xVLLk8iqPewc2Zah
Lsz8j29qq2bcPBQJracnNTiBc4ZJor5xWtTDGndh8cC6Kua9bQncu5/9IUPULQ1oXeUBXlzg
C0Oo+CtkDu+HsI8Ce7+CNfb5QhJ9Tye8/lmSnNaK9cr5zrZwUuY+bn18H7OPMqlRJqReB2lZ
pJgNOrLCsV/EmVuACtopEtNgpjBzD/TYqIp+Q+MJOrS8lZvIz4DIJUET+yZ0qcmSy/8mBh9S
26h0h+8m0kBguJIwUdVI5jv+xjjYPlvaHrc8cr9KIPY8ncOJN0/LzZIf6HFEKURXXzxY+ndh
ChJ7per42iQfvxHx/12SEev0eq4bETYefo5EfTANQ/fE7IzxLZLflNhmbFFamWfqiqirCQZt
iCLwZesCkrddtCa5mcCMVckuV1BEIxTAQgDyu5Lxgcxb8/cQzFCbaXlX/2nSmN/DUEeCRS0k
wODyhSZpe5/KNT2qpI+1cbrxMmL+d5nINUuydz1FmbWxwx5s2tCcUbAQEpvoeS2ehT8vIBBw
rcZSzEejaY2ih2+HrfG7FwOheidUzKCtRDkfnhZjFyFeHdv/DzjCTbtAouK4Q+bVHUA3ZurH
ArPHBgkwOCCjaHES7EJ7dhXbjOfYZGjoqgL5haRr9y8olYFjJeZSLOxLTfRS5wmkEQVkdsv9
1fI04XpkuK5LGvbeI6bxyQaYfumf+hDHAEQN80iN+mg5VFmepEJgMmRmAGbRQE8FVIZu1/Ic
BqmB/CMfCCmjG6EfYQ1JCvOObc4DWXExxszLLQbyGYxpVMy6+GzPqHPhtU1pmGufyN9p0Z6B
efE95ZVECqIg/9U5Mzfd4L4ldcXYs8NGQr7tslP0C7j2Qv/olSOHVmqbSgoGhMzjBq9xbdiM
bjgU2oXDpHPkalEZdRomHTq/fTdCjsO5SesRb+5eE+O4uIbuu6d/YZDW
`protect key_keyowner= "Synplicity", key_keyname= "SYNP05_001"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
XcmkvUBwCN+ZIhO9GRz8NZ0nyInROk4wu4SViRe15cN2zOjJHaKQC2L2yRhR0x5X2B2hfQk3
VkIiZY82mRYIKyW2WzqVF97L1CIovnp1AHhPfce5wapbf/xF9eZybrdOvQM7j1hsTj/24eT+
2lvyMnL0F6pr7BMWejmJC+DRJY7ticIENZ9LMfvQqlI2Eie6WaXGUYt4stB/fr8HkGKa4M1H
/zyhgNKXFO4p7xNJZty/d7NBt1YtVDlBJTM/hpISWT2DpPOdWUQhC7I4ZmpAkAIaNPBjkpX9
14NYNfnRLUhL2N5+XPkX2LDRY1hFA+hCeqbwdZcA/3FfG2HU/6Aedg==
`protect key_keyowner= "Xilinx", key_keyname= "xilinxt_2019_02"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
UWDiGU5jVjjA2ruMHDPpROQlal+Hk6iDPm/lhiEPvzXcwhQuK61yEDJWLZPv0Yr8Ms/peL0Z
uo6Na52i7RIOwvU4s5K0cS8BoaoNoJGjhFAiqHlzs5p5/KtrND4Abf0c43iE46RpC0G29oIp
sh5HKhdO8sgOstS0fU6SzW+LZ3nrwoWtnHy/q5J+bUi6v4JX4ZLr3PC8d06WkQhMLn08hYQX
U/JJsZUYzVrQg5iCPY2g+YeQkKw/aWTNkw/uz6niSEcquW4jhHXuJI4/Vth3OHszmxjBP8De
OJPKe+JWG//Bg5fcThArEpRuNLVQeJGZolwVK/q/MDJqVWnG9JT9mw==
`protect key_keyowner= "Xilinx", key_keyname= "xilinxt_2020_08"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
Xmq6FYh31BxnlPnJQZqsboYQcTcn/vyi51c7mOVvClgfj+iunp7c36m35JfKolGPXRkNrl5h
mAxU+hCIp6fRW2eCsXAql2OLeR9hmUxd/CHuW62lwjQcrFVENEFa+2YV6E2ymeOq9vsXKTEp
dQX0Ldq4n4BPQajQtA7DOrzuGQRe6A0Louk3Kb/XQI3uri8fj2qbLFxb/h+0++dLl2hLmorL
vIAhGj8D9I52gZgSj/Y58jQEdpiZXON5uQu8sm2aZXtl1hwAobSQClEZ9zee+0LJWbKMNFYT
WJo5JQyzOx7d5P8jpa3Jk0RkhBEhQyrGD3jyzTzlPEHNgRcf7G/vMQ==
`protect key_keyowner= "Xilinx", key_keyname= "xilinxt_2021_01"
`protect key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 72, bytes= 256)
`protect key_block
jXjWnzXKiTk3YAbvpNMxoeAmlkVnTN4nMU2yUnzk2ePcxe7dmEqKx763SWMWVk7NDzOHnW//
ipFLy3b//0zcm0GqA/o1kg0KTSqp7vbcfSMcjq/tfvZB/kqo/dXOX+yeaw7A690I7HvO3/FY
TVPyCyyxPNGn3GfqayH3AQC2zSYdS2tzgQ37GD8vJwLgUx7eePbrZcXqOOQeMDDVOVcBIiDs
Ua7vbcHhLX1MRR1juBIchdZdpz8DUv0YIL64L2qDCD+rX5Phh4t+dxpZ6PXaTu42DW6LmMkC
c3MeY8ekHU2qrCVjFcTyk+Pko6e3Pv+KmEstJ+x894g9vRRttXo+JQ==
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 72, bytes= 25216)
`protect data_block
wiKSMOmn4lY22gqXf26/c0xveTEmy0ZW9vemEjvs7RWLm+HV4K5HgOGt5W3rb//jDNyf2tbj
eWPMWq8Tx/C9MbjEKk1L/Ip7TRrxCPuTsyMLsH7NANExS3hvFmZK5mYpw1eNCs0VMN38Q/Bx
gNsN9AuMfPO9WNtHO516ZoHPe8E/ifyELL8SWvzaI2SDMiHy7EpxhRztVFL5/43dXZWY40Wh
3hMVYY7dvuGFdak4oT9QfdxS3ncyiYBoyooDXgMx6Jx6uY9eVN20FDSNTCqODv4av7jhC1Vn
QTUy22KOKpaKxIt2UStC1/S+PZ1CS6Z1b4CBnkqvaXEfCHEyJgjcKEZV2ZH6OcmWCxtzS2WL
OvgZRKkqvM39rkBbgik5NOHdUr7a3hYC++4cfqsesJvXr3/nvRicW7t2l+x0CII5HAIu8AyH
Nk1oSFSofLh8SAQYh5dW1f+2GYhOLgIf/2EMtMhbRp3shJRi2TMLFwCL4FKjBbUjRnzicYRS
xIXhZNNmLhtdfBd8VjvNEBrclPENqTmlmEiXp/NnWYKew+9Tk4o3sKZyW8d/vAsSPNdIe03m
DHGasuHGG9JEdcGlpoYQPPWnBdzN9vsOZUsnyF5RQ6+7UOTftlDw4cJROQbr44eR8p51mQOR
REPs6BlgHWNj2u3Nky+/WOvM/ombHOxObd8L/aB/5TUC/UiC/5jh5DONzcwpUbRWD8tF2wZm
BoSoX3cdzySOWGDzP8wNCtuiJdOVmtfwzC4mbpd+osrQmMw6uwRSHnW58EVq3CJhzS37WxrA
3YSyHChNcGb7tDoO+XCruANhrfRFrFDwXRfN9fL5qM5MwRlFEdOlipktxqIwDA3+mRuumn6X
2fArpzeAH12H5k6t0MO3uXUvoiJBs+aEwVrCHAgqA8cIPEFzqAEubdOxPsnm2F+67+3M3C21
z3L2G+t72zYEQlRCqxtND4PGgfFtUIlvIoJG0QkFBzLzEufvxuD+JSLM39HVIuTaddu+CKNO
zdQzHxU56GL89/eJGZMbSDHy8l3xTLBR1nNH2kswslL8rDI3eGr+2CHDMRXMMxUOMxpn4apg
RXvVSwOsfklXe2GnboZQAQZfgGAe9J6aNVx3BDQDk/ucmd7Mb3i6J10Gu7spdS7Yzd2VDMdN
9kNbnoxMWVjcAezRDGJWueXt6eXykXNULp17dSQ7J8v7ZoOw/nnUNiFfhWc8jRdLORacez4T
4JVVioSED1JDANEX3zkD10rCgLak1OO7z4SON4fx+qE9T3CiP3unYvOpaX7CO91zCXkOZRk7
g872tB69WorGzfUNpje5npbKbApSqLcxPhPs9otlDoKkdWohyD7QqTGzkTvcfxbj6HlMMFca
EFxSYGX9fwzeJCuUFxBxmp2mBlzQD9OE2jQ5XdYlh3voA0Z5NGogyNq7Q/RWNxkbiFgPT1Tv
fZQ5s/h0mXluaJZ68nLtx3I2l+eAaj19o0bGDO938OasaWUbKWcED3is0CAbihBrfIeb8nFr
6EDhJSsFIrI/GMnxSByI+QpDmfR7+j5hP9PMfHlNUq6Kc1zkNKJxcq9uFbBW0NqVp11HF/ai
RViP5Z1UobVbnymDRKfCMuZKTxmA7t8QdhIHr/RqSCC3x2CdwmI/gNy0qAb6UfydFcxYvB0V
KD99b2W5BfVqCvLbILj2/I1cM6e5iecKdFxzDUNgb+NWxSpzGplhLstW7R/A0Mt2hUSJ5Jj/
FxtifxjoAuiUThfhIiajYpBtnnXIayTEnDFYi9WwpE8PDMx7fqhB2EEKo9XRS8j8WtyFROWj
fMNLcPGSa7xOAafz483lGd7/gKFRZGpo7f/aU+R0kwdAffavH7A768vkVGIzOc0JMoV4Yihb
Erkub1QQqNzSJSomLbiDPmuGz3aOJaash/BgBdLVilhVDx/RjW9zHRUUcW3tPRoGDznaHFjH
4RQny/qCv8HLyGefY2w7X2rNYjEJhLLKBb1f3YojnuFJSs9JsMfTvIpqVvWayJXP1cBzBJsN
bD0X0F8S7TvtaK/NJdlLss+6MkAwDXKZ0z5BEcf+G2/9rHlObt47vjLyZ9lWT5mo5JN/bKrt
/KU5eraL2FW31j9bOPSicQY06XX5DRhjeNiy+cdIZqxzHDT5OkRd15ZFaMtA549YwKXdECwS
jFV80iHu6KNof/ulgf4sr5eGSlO7PWng1uL+vkUFeQlI+iWsMnRUAdrxBekIIJVfFPe1Sr26
JIq75Uj48vpCx6sNUpIKKjG+llbnfsjMwRUu1Nh6beIuuwj2T1YqPWlVDVkoJlcEq4fwt4yj
MXlhHlC9r6LmiJtgl5O0sLHdv+MTPzRH+9gSGRGnuGgOJVJvGRfLgglxVpz7F2Poq08T08rA
6CDHFTmYuPMdGMuaxlQLw0rVd3K2e25xHQpgy0HnNfSpk8AaP8shtlT4FxfTWDXy7D1PJRzc
jrCF9avKnWMSk0ciKzkLHAmVm+3VH+SbqZ/oRgL4eJqHt2U9uI1yo3emDwDYpsQGVLRMd5UU
VvVAXWZXdlvNmRjTSpPaLPBCUvroRBiBMTz0obiNZzACctSLc5ZNDZzkjUWX1io58QOvfd3B
55WrujOL+N89RIO3qQBGWhMYof8i/OMs6zvb3VIkyuk1vAQjkNjdaff9YOveP53nWl1zTUDZ
tRAaHiiuj4dIm4Ce5m0DgKlzCvBoswAOXsba5SHg32g705XEIK+uokGT0SwBBs4s29wLyVs7
bpWEdVOjxQ6EMGOadr/uWxFBhG6n7DnQAo8bS+hOdxe37iPrOBcvheKEr7ZCvpihvwh/NvoS
6k9P+xEnK+NQOiZP/d6kQgtZPCT0EUfHNGgidMFeT5dpRbXWoPGXhXxTza9Pvqd501f6iSn8
gdAuyCa1OsEv1fotJutSRf6iiy2vN6Zd+v5r4w44fkawHzCT/43nxASBjpBwTKempl3WnnZF
kx6Ggu4bIp1hXbqCtkprX0KgifVPEaCuuEwN3kx9/KK221bmniMHmfcnej17q32zijpntFVq
BagscXyxRyglPGdR7ZWn42Ytc6jWGmbtRrxnC37fGnvveDTOPmBwYXqyLR9Pe4vNUl9vYXk9
kzGvOM9vT2Lb1dUsOFCvb/1vt8nUwXLZvplbTotgusgW2DOxFAWPgsSRMkg7y8q9HFYyfT7n
c6uaeRZrc9XdHDLAu5jSXSWKrUtkcY8lc50Xnf5k8hAFwBls+V3qjBsbOniNGFgugbD5pLty
2ojC1Gh4KfExS7mwyoK17fVx+XJAlmUtahJVdi1y7GiP4I/qBBWyNZfDFUWV1BlRBmx7eWbD
FCCmzuI6G+iHYHn8k6crPfWSVXdL/WeQuOW0ZeuQU8/nlQyiI0o1/62WgKuulUb5ab4Wg/j+
UffQiIHEs+kdKg0wPI6XekK4n9+Y/e5ijAubo2E5abXRi1UhWXRqlq80DdPEduKO0nM4xX0z
pexNg8JzhJgevg/+/9VNErh7+qnOGpbdjBFtVJIUp9hWwXQKk/33XAl+nuNKqAzAIYbhE3nv
4m/31vAPkRuZYNXncjFDsfWbJfu7HMvhpIQatp+U14sncX0k6v0RBXvSU70kgy5seEmokRWf
VkVVUaHWkxS5cNka4YFEV+yzncqmjtSYDO2MCiqPiZt5zxXy7tH5Lu0v6Tsc0y722Qe4RPHW
bkkGY492WcSuPO26rbtJqa+XJJi/6aB1zwGwDfMOeGmvuQJ086NCgvsuRY3CzZFqeDq1frrz
t7XEW777dEQkyNGc+WKgiKASNojrrRKA/ronpIcdh5o5dqCiCW3NmDuoo9wnKocIxE8whUug
Kc6pf5Hf7xig7C9pfQE4mBgP4gNgXnPcPFaW8/QRaD/MNEj7cuDqPrIrGr5lncJTYLcS70qY
cJOdo6NnWorI9NCRx4hTd5yTEtfj+o/ec6Na5th/0NRadL21tFeeSPGgHu87yR9BDJ8Ko4Jo
pILAZaaMCWGD617aDCpkTGvoCAmEPti9L2IdQ1mkn35M69vqzpjpIf6L/bakbs1/fcsigSaP
oR9oQI62cWy2VbnTZUXx0uZhfm2PNuOJJNVHmlqf3R8PW1uITac+x9EzKZ1nutbpN1tf/Uq6
L0rxSRBVexTVDASFXshqpibczSzJVDYth2gKwFFBRgMtqjhX5UFRfI62QIeNmCEReWzhuLaf
ZJKGmNsZWi+smc3uew4gUfldspkyzh+KwVNUwX/ZeHWee4SvtXpFcWAkYCchaklR0tR32pM4
GiZYyHH1yR1dsNwKzwetCFbJ2a7HeCgD7h6WUi2yP5gqSWb01nCu60+RHtwlFuSb8/zr41N/
7SMF2yRGjqUENuK1lMgN585c5D2XoUmp9XDoEA6TL+2jK2qh7ij67c2jDHv0fAlAsVXGmziz
ANpDxS5J6cys6lbmM8FHe9HevAIjmcbLsE6lna6l6k74tztMmM2zk2R268FsRPoeuWHmwdQF
NsZpxzPQDJFpZcPND0eGLvqJRivxWzhDAGvXZ21hbUcIbWYMjMQLj4ZJeaqFIhdvbSLdy2/i
aAMSte4/5qQNPo+I5W4nR/pc0Aa5uX5hNAKAs32zXTvWPxJdtPReXEOS+Fh/fqdRrHGHLt7x
eC7MoDso3je7DrpIhqKhjOHIHrWRHg5MeNzmevrk9LvV6M5piV5YpNlBGDT15AqhpOY1lB8E
MAJ6msKjp1eImd7bnR1OTFwHFEsSJcZ00zyQVdVxjPcAQbGZ4qIYWriIM9p3Y+wX1RGAd/OX
ASUtdXt9hDkn61aXraHn+h3fT5GiO3u75ZNeZcVP24r8rslBs15RngGKdc4a+HYRMZi4G9dv
D8lYyvkBJCMNG2OMTCt2dNsThkV3xy+XuWnh5/cnnPcQo1EIzux8ArdZIFN4n1OStFwkup+q
LnbXeHuWnlHl6091RTPWcQOp6Fo/MUiRi0VwcNl+X6w+JeVEi84/yzXiETyHq4f5zW3RLRZK
9nhWAU3y4pASzi5IXxO7LYJUYP8k6mk9/2DirjdUKwsYj3hOq8bbGJjUGjTgzwudA4VHt5Hr
Dm2bcV1SY/HrVw40001tysr4aKxrJNhCxXr4KiTj4o+mWZ4aq5CBUIEumFbKtKjgROOrODDy
tHvdYiNUyFIvja852yJypZxEueyt8ggwAJmIFmZbAo0ODjT9e+5VzgnL6Jqa9tZsaKuyFIdJ
ujXIpeUf2OTT+5KSRZxuMZUpJIA/jAH14HzyN92jHwm8bns1l7paNsi0i0HtVhgNidcJJat3
kV13DFOb1fvHkDxILl+RvyuvmmrW8WAq6RXDEP1ffetD86xsiRsHGRSV04M9vh+4RRSMDaVh
dwViqaMLMj+3IgJFxEfvpb80iKA3VywraE5eF81rI+zF3UBibH0WerKUSe0Tb9dF9TydyLn5
UEwPqx0SauUAM8VjUtFb2m3Ay0aJOpgOFY5Js8eE0KojAYn2l22sC6cwc4mAsK7MhvZ4iU+n
SXHFU1PiAjOzcT2nCKp/RrPKxDkUyOFACFfE2PgNYX8vmkBtvgSM7ztaGccs+v+lBLdCmwHU
QmNXkYFgiHCvrae38zNXULqk6MKgzidwoyNt1DKe6VFHzWRJFsKIsuqJi361p3SxtaCaf8ET
E5qZ5sUfMySnHqSlKZ2OOGfmfyRrh9s1eCR4pVZeCc2A++nesl3AD1VNDSWco5E2yoPC0VcJ
LbsqMKybeDuyMa+KWuSlIwcrsowxS8oIXfAGb6ToXHSBAiGCLQWXuv9nG8bEUJHzyeneEptf
RbFZg7KSKbnYBKYtKzts+Djsr35+0vRFWxPOChKg67t/Fe+1ODnTNXcneAQhNPxZbM59L+Hu
4HJvRqWawKPnN1VeXCZIpzghUL/rswduHw1s44ndaYfRxqTcaerxtgsJ4Mvrnj2e9XImIxXN
m72pNl1dRbXCRLqLBGD1ljq6yS5YVCumjqM3DJBCtzNwp/9tyMQweXPN2BbkFHOvsWQsjAq7
tRUUAmO0iWyqMxB/t0euBL4bJGC/+sJDrvOf6Dws9/RE2ZeHht//87T4lNJ52PpPq9jdHhka
AocxULZGiyJgf//EogXevWxPnA3quIrcY0EwrBbwZAMYbFASEOZVeJ595ZUzKjRxJ4X7K+Q9
WM8/qv2ejEaflheJqRW37M+qL6OMrlGRPfawUb0zg6RzY3eDLvow2uzwryBf/uO/Zy0kSBCK
B8q+VrsqF4JrgoH5DFWB+d60/G2slVavhpxGoMysqGwc7FRECL1pXcQ2Wpb4f550MEJ3ZstE
hwtaACPUL6MSRFWfroi45SJfSHsrOfmXDSUlhZYVfZckZRlR5otudghRglb13SCtTH3fAZ2+
mBHzc98TKJPsiF31I84pSTD91bFliUWuH4zXSmhpuzKEbl8GGeTZoPrt4ZarpKaY24yJInCJ
5cIjUB9UNR11MdtjEbtbXKHpAXn60bPM30XE7Z3wbxLeiNc5ssAYkbkCnRJwnfnS01N5VQpr
F/Y07e5hrruKGFYmDmMwNw5pdOInXPTx3UEeSu41ElHUtrtzcKaUj8N16TvQ6oISOF9mIR7O
WNo92rQXQV9zZ7S6UoK/fPUg2VROoofkvd+mMJoriCz3r2ce0ADJdQvdQUs48i4eA1i8sviq
JdSHh13MRTGXKMKjxbKNnwIf4lpb0QqdsyE7Sp5sbg0ZSItJsFQgQS7lJQZ/tO4TZzQnU47O
Qdtlo7u+jdd+4EvHvCOkMrWEIjrrMFKcwSuxDW9mJkNNw6U/1pHX4jgkuRCIpOtLpT/hM6Ie
7BVB57OMTTpP0dZRkHKJ92P0t1dbQLVKAoJu1VitqwjP3PiJIs/e6fMFbiP6WcQRPoJqPpQp
RGKpq2F8GCM1iDwLqga+kEWbSY10f5Q1z+HOz6mr+Nj0jscH00QvUq5j9qNINw1cWI0vfDcr
ZDGV0TopatBPc29wpuWRH9yGWf+7OEmHz2G/eGkPe2GUYF2nHo4842B7YKX9hmLz4W5cn3Xw
C1I0VWZDV8GUp8YDZn4WCn8ZjzUHK3Jwtk2qCa7P/iIaccKhWJzrvU21w72BDsYpqJ7Pxds5
5ISYm1XayKIO6EIkJDUdm0kTajZIvFES8o31nYiTDZk2VmWIrnm+3I0yxnogf+FU6FP5081e
RfDQFkw4OBz6ltdKuBkPjaWiM0xItBrpbr7IeDu6EkQGCp+8fbu5Uvdfdb54GuyvGV5C/gjN
z/RsLjM0JBTVQyluS87HI7+M+xtHH0gYTz3R+Y9ZFagToHsByif3KSlJ0DmHwkyIvBr6ddGU
Rx9jzCkN+QWH7u/Ee4CWDKnjZbI7bMKnDhR8CwuxQvV6uZy4tEFFJpC4UYnHaGkgvFw1OpSw
S7ZPzZkTHEgYOiKha+n8YEH3tvj9DAZxlKcMWBcNkMFozkBMi6mBT0dK44Tl2uU09yPsDX50
Q4P8a4L8bCJXZnMAbCBuQZjqCeAGTXjA/VlGMJV/ZmGexy1QSyyWz1rhIDwr6mVgfFN16Z2/
ahdeNAdplT4ur9TvXbOOlwZw/OV3u6FCkWtW5z9GN0diMMh55cS3kLNOuBe/Aqhz3qTd0MsI
c7u9uYiH88f7991CEWd0b9GoFCUfNvorq9qQ0lIa3v9jF0cnVIViS8fEj2Vth2kw5MSGyShw
/tmb8AJfPHq8gDGEsbaeCrGMCsEpQX79CH6ac2c5/FdBEgCfFOMqs2oMZ4ZVJtUX8xUNvAm3
yHL81lT5/S/j0K7KHgEM//LMXueSoLj25jy6oLMkcWBtCarf6LERGcW+VIg/CN+IbyTngTHN
0+VoDS16XKyzgtpydsrOK7NYpiSNxxzCpRxWvS6gM1QED6U32INE1U4lQK3CLUWIQmjzw953
g6iHmB3BcoNG5vyeR2T7MoqJLhhUXBuy94CErh8LcoF1NVNfYYHAa2FrZS7EEPrZ/QVSCNK4
n7pyxtP7SrW3K8/8Yi+IphJRcTq1CUVspFFQzr7OkTsm2sa4mNjsa9OYBUJcaJSdkz12wChK
vRhiyP0ftE/rP6WsMA6brd6EBb5pWxfR6xwCywmpSDw7c3kEwbY2l52J4kg5llqYueQdCYqd
yavqsol3DfdH6faQbSUxknmFUtT/yTC0czYapcuGx7/oXhjOi18yY1+ThE4f/BpR/a6VTWNE
v8cDgbJ8xtitzJ9JMHByjL9l2jrCW7XOBjjmBYXgPFZgfIcv0g/RPgTVU0WpNSZicNrcnEDa
PQ1ftY6Gqk5wuf3ySFF3ljz31OkLS0FiDkN24JbH02xXeZK7xc6LCTCNMlA+GA90LWf0xQgl
o96kNQH/JgduIjmg0ipLEIiJC3ls/fK11s+81YMgV8SM/WPXhC3pl6Oykukilom4kNTJh3bF
GjPBkyWmGB7helclmmr4OGhak45FqOo43z03J21E9stH5FP1lQeZgOPWwMkBjla33OU9rQG7
aODM91JuDsGShyK4CJGmSU/ZO//l4dpiIQcv4sAmSQ6LThRmCOfx3MbyixAGC2bbJq2QJ1pz
4rICuk8Dx3UQiKGy91Mf10T/5iHhyBww41WD8RTpfMezCSG5I1MvlZsqsM++2H87Vxdd/hBR
kw/mPWXLu/GD4PBEnkKCT20y/JS91RyecklpPzGlJZ03EaGdoLLfj36FqF3fsv59cU1mdadJ
xtp1v9OIyuvCQXUoywT4xVdrUcSx+hxYWCxXVB/rEorC515ydYC0Vj2ZuB4TlijX6NJecwj/
BgyOBr6xr5lusjLPBa0xHAUH3VgqaKhO64A22ewmrx4Z4Ne/uQGql5dZm8p+l8bkeVZ8yFty
zlSnySX0NUBWSCVWea3MknJNFRko9bsurfNDEWNsV2//9zPZiDzr4CwMnFMjFSYxSLvhelfh
zjnvT2nCkH3fkuofbnDQ+tNgrR3KldFYODTf1f6X+0kKphXRzfK36tDQ4Ug1Yhnwo6oB9abF
qmNVcBpXTtFq4Rv/n9e1iVO0mNDSqFySrJ7Wyrv0qt3j+eyDxotQFqsMXhaGzKeWKyMn6gFU
xDkCWvcBULJYlEP0K2gIXQSargzCju0DoQPDVikzCYq439H1/GIEgqNmGoaga+4KCzLdjG8c
DUHCdDsi9ds8wmRPTwszb39av0aZ0EqHCyJXltKqfSgMc979FfIjjXgJocNaQF0Bz0FwdnjC
VtBJA5r2drBHyvnY5g7GdDHGyr1XlMc2oo41G0Peu3jdNtmfrzzz859tZS02paehcjh1zOAI
TpqYjqHp4OnuV8mcWQXvoSm4ySD0uFXCe/YpppK+977RAO7TpQwHNKzH5armoKjXMEXWQ4A1
9PdbF08WmZC/Byekqcwn6GGavV45jejhPFvjXMcpkcDEURcxEg5vbtDDEmEcEABm+Jyl9wav
XFVgzF6GXrkJZ3KKSKsYLgj8u5r2xlpuFjhj1f8PEMg0uXLN1IlX6PNwZJhSOqG57dcsGt0I
9eVD0W9oHM6lsYRK+VkdeDpHLJoMyLJqVWBdzbgJRWZHxILnvbqyaZFv+0nMGHeP0NHMCbJk
e10tFvyMJIDSOhAtmBtmN9jDMB6oOSF275ds8l4TlAmAVmGj+q3oBuvrNJjRtUI/b5O2SYNR
Vxtex/SURWp2usBAuxCj2dzB/ecLN6VcBgMuVdfKfOVg3f19/Sh53bkgppkvY8mR5Ob97EfS
Lk2kKbOTLouroahejo5aIlIKwqIux4mIOhNrIczTHVzsKppNJees+p6F5ZSphLnkBbmtCCgf
FyK0pwVwpH0SzIYWxbhe3PYN/Nyx11V91oxzXMbfN4ZV8W6V0XpGydIg3ZquCDPQqFO2Hqv+
RGpq/nLV47zk5cooMOYQCd3EHMfooVCtIAFV/v/hi9GFOSOX18FXhk6ipIKll2qz/K4N371R
Ahn8bqTNNg7pHQ+SGJahibm0xkDb7mEGls3ByIcM2L08UwkDkdMv1yhYXb72bmFBG2hBDOmL
GESo7x0EX4Cn9N3rengLX+ndjBvSr6TI+VACsVc/3wiwjXOZtf3TXCH7etIhMOsat6NIAcrG
IiHXE5WzoCyPxZ79nVxBZD401Hg+6GV3FvfWlPLUNXmePNG189JBeeQB2A+dbEobRvXac8pT
PXV2O+Z6X7Q/HebLOV1Omepn4xecv0BHI7mvdm9gHkNf8RdeGdTJ/++z9dJUzNEgLBiAxBOU
DiAxGudHucbRvMPPEwGJGN/yiMWxxCplt5P85bNXGkAn4FFGUVCpklbsEofEV1vysW4fuvmV
AHQjbR/yNNih5uqCEt2aBuf1cJuKthj58n4wlgBMx09zlM1N0lX4AmaPR5Ch9tG6k54mTL0L
ikd4SGlzkUStBXrCkob3EjRAwZsTc6vZKO4bOWoZ1ckKcPQmhkuIP63mvX3zV7un+H/mvPGn
enSYJUh4o14GVTVkIlkxGIBviYOa2wbyhbi/AO3H+1vH3mc2Gj90U8dwU8/GlkM75h2IQ1To
1mGhArmSWQs9WFeEEooaq5VF+Jc5ExeBgX7ba+c2Cm0T9GuwJTAdwqgN1v/vMpkm7u1z2evl
LW8iramq17HOme42f+n4nZ87MBpPt3Mi1NIhU/QmRPAoJdYaApIms8AOlu+MD0fVmCTC2/P/
MtHh+dljxrnw+b8p+UA/D5AxTw9Wa7X0v0xixXiElWMGd9EhM5ZNZ7xbXOxwIBAMBr9cx0DU
yKJMdwnqxQ9F6ixMq/BWjbhW5Ljlmsy3PKawzOeQDwPOT7EnTADps+dUiQNOYPdlVdOTREZh
5/R9m4INTFpF5Jro8xkOlC+GBsllVLLzXNzPh8xBiI43aVbSUJUmQalDjNYhSXSdlOT4JScU
H/uAdr9ozBKsT9X3J3bUFbN0eNrNwkZ9B8gwBAsyS/wfNUW03Rjx/FsiWwMZ70PJs4JOoTZv
5tLHjNOfYyflBQW4dv6umBt933cEbha+ptOkB5RMLkf5bbg5SG/C4kHU6/4XXTxJNBDseWuA
yxwHmdUHp1900EPFH3VHl71kwVhBIUNHYPpfapev06dUjh12nmesT+X+N0RlYby+qq1AczuA
IGWw6W2K/GyCnWvMiK1EXbDitrLc9bl0v/Lty+vVR6CxYZF3lpGiujpKTlcS/tEFPrkTjfmC
k18O4/U1u8oNl0v3YErSQzfhCKL2ZxcYyEfSns62qDMwTE+H/juLFYwgIAeRRkx6JfAzWDCZ
5L+L7JE4vcJ+Mkw0hKtaNW1iXa6dTKZ6+Wn8TcP/h8QhIqpzMJXYPGpyHUL5k/FldrNqXvNb
YTD9y7DUmh/ZdTE7eEy3da5LhWRi/vqZloF2XU9jLieL26zg0TB29o5+G1eDw9EwlOlxufzn
QZNOvsVmeacLacE9f/teOcx5mevbf0KHYIusmNr10jKpipjAOFBBIMAUSxJsC2PTH1ABSuSK
wTl/dssq/V5V2V3nNG3k2RcbKZrl3au5giP5bNUxR0TUWFJUkcSmvsKRWXuwJpC3rf0JAQLa
2Q4O5lKumGd8AfTaXxwmtUsZysnEp+Tql1yp7nq1Cx9NdlY07lmVj7F81Gbd7TCFFuo3eUnT
Na2bx9/SeP2dyfU5ny6SKWdfHXVvAKdjPxHdz29y25fP79ZeBowcNA25gxvDepB82VSsCxTS
AD/6YR11cfjuJZrPwkOZEAP/AnidQa7L5o6gid7imlTalASWmoGgDI5Aem4mF5FPliHHicua
vFno90yo09IC9ozDCRuMpM5aKBhRnifGlqXlYLm3Y8FYG0LWIKnEN/FH/0EGO5Y12TscTEr5
Ct1zaWVNTAaXq3n+keunJ/snbBr8xmghUZ+lkeqO1Ya25ola9sejLIglwmdX79pQChDuAQui
AxW6j7QfS1I9LBdkFIayY8klWPx4acyXsRWI/4EwQ8FhryOwBCeEpxgdVap9DcoNcKJkRDCB
WAMfrTUVujBYZ/gBfZGtIEbxe6H1HntgE8eOopC4M8dYdO6gIK9+G/GtVG/NiCX0aOtS5953
7NEU1NmYYNxOlfrbaAtyBACzX//YTBJNLZqLw2w+TVsgNkV3lEzjvW8a2hXVuXGGlfPm5o29
b0oUBa/S6xQtnk6RP/jieGvskaQil4s0/YFhl3jWl2l5jAU6+KHICRjjy0BOmIdXRt0a80jw
HcFk6e+F2WyXGIYNpmW1Y8RfQmTXqP7mHcBeA0CERcFJpHp6zvO6y1VrKF9Dj8uuOye2HPVI
NQGGSVtISfngGUFfT4sN7IVecbGROF3+ASMD3AvN+ZdnS3gMhW9DT9nHbkS5bo3rzHD6MlI/
CsfD0bXBQk8NLHnhEtrmjoHvGzzH8sfafuQqfXu1JWASnhCKLiGm0Jn153oT614WlC60TirI
IT0irMu5VN2+wB7VV+YpkohCVJwXMScQZ7fQpFqE4TGBG3f/47/7QK5ReF1h8vOf05upHlEn
X654InENxAs4WEuwifNYpy8ojOimWjk/sKQ3JPPiPTzEjMGD0fbJ5Jhvv4gu85cL/HoxvHM1
2x/2Z382ghca714+CBJxWTHVwi4RtuOAkTFaCMXv7+hvsUKRRjsJ5QOXqGBWr2DCx7Z7MWyQ
DLIUxEpCtiI3VBq9Gz9/G5spztr1SA1nQKEKdDp1QFjRe3F2qfLGWNMtakWGH+LEZ41dm05M
JW4jlTX52YFA5QPntSzhkYv32kzRK3QKMQe8XdJ0xDsYLomVuNACUdb0cHP5/ZTCOf1fpFKV
ibmsrnKtDLoRviXV9JuZDRZxUQYUWuedL1c+v8qilRePT8WoORIILIUZH8NCzFka/b6UMzS8
WMSc0PpBxJmuWSrwVdhxo4Net71wbn7G5+xVjnngPtrc6H1eDwYS77DAkIHz+/XM2aZJa/wM
QkCo4YIQ01xSx9A3uu/gJ/rt3Ed6jaSHqGPU1x/lRvu/2ToOF3i27JGDR61V603lhXKvDKkM
Ktwp99KXKiZIMGJl/vl0g5US04zyQg1JnxF5lbrRLa0tSdF81HQRhXPplcETTej5Y9PTY2yF
+l4Cq2/cd5anQ1iJqrp3wFl+dJYoRvibkzLZRGDioCPBbQ9wjDj5mRElVUkBZ9aFIAQhknuO
UhgvsoE1Zzy8teGfodYEzMfA2JhAbMSJHKWSbShpzpuPfYrst65FDLKkMqDMeYObiLfea+14
SU94bPbPNYAAse4GaWShI4GGHBH905mdDtjLIBdxJAIoH1WNvlIMQEC9YU77Fy1sDgI4Yw/Q
CgKS+Vpbv+xwX0oklhm0g32hCV1LE3WsQmQviMplGBuia3pf5BxmZ45UT/FoQ1gZuHCMw8ZX
AEU36u0dxqMUNXQWnQ2abWLm+zTx0dDiPw4BXbiqCCr7VN0tPWj4F70Tv7Xq1J68MY6LC+Y8
ceBav8HoCGdK15v5WknSPF8u5IynFAzCRpLZVMSPGil+wReZkwchBO1N7fNUW8Ys5Uruv0FY
x5rgnc9Lj8eLczs2zuPJ98ErCJkAMkInJ7m208+u60D+wc5cwgBhl9YAn3FcbmPXM95TbjRO
BQ/7DyNy24Y9YLZrV54ltAQyjpnxaSacup53x2Hna5HCfWnY7udHzSNKRJKGxzFsCGpT6PkP
Vg/PVWmnbY/nTDCq2TitdS5Rx8rxw6bPaxfWhkuePdsmLQVlny2ynx2Jf6FHbAqoYlkqCD6L
oCDu1cwixRd5AVDvKtaxmHjuFp3ZVJzOEjd2ZDdUdDmLqwqWOQGEhBNxm4gJPt173AlMgKNT
vuWBCYxehWuIdNfMupjS8pR/ugE12706kSzXtK9XQmyqzYnmdacJVk3PERxPx6LKe8DQJGjD
zBa72nkqbaSfXUGkOvd0onng4zuEIzxrZUDM+znpN9grIRc8HxelvHimGJxpiuuiGprlfuo6
1QKu2Av1IhFPRxgvGu16Fg5I1RhoVfA/py5iSlZZNBrHLEUSae97DotGnftL/Nr/1DjFm3+z
sYnQYvkBSPwHNasjKPfOSOVnIsc8Eodsfswa9qZj5/3YUW1svGk0/fu8WB2L/yyK6UPYf9Tk
U8GDAvejGXppAW+Hsl8b/tBkxpLYeJQfkhJ9sYlIFqugZ20/wQpPG6w9nfOBixIJ2DssHHv0
txLx8FXlH6yp6Fd6Pb/DEtP9+ByXsYOMnE+/FZBEkmlD/5KQv7DrJCr6twSqs0BIGQE/sKlW
szyoiXzlmpje+yg1yNX2ZXTxblKvvClcpN7aA3tUZlknG6gO0hIlL4K+Vx50oEDuEVXbAaRw
XT4ckVtZmMyYJFvFZrYiUpOBfDldyYi19B9RrBV3YxEVTNcEaYn8HIXJq/vSx8p9IhZDOKOD
ijRUWEUN/yDffmg2iz9uKUGamwEn2lRwjAqtmRdUPQeXzLGM+7TRoVFcGMNjlwur4VLgAY6Q
KO69jfQIzN+5xYBj9J4ud+LiOaMxXeMORD7N/9oRs3Xzq/22p0G8ZBHy23jLArMNrddwb5LC
dy7OoU7wDCuBrZR3EGHWYxqovdJvjp7gkkASbfY2h4N986Nl+I1TiypQ2nJpRgQhlaZsdkhX
Mq1iOTi2FdnL6cR+DH03kotxmRJlj89oAqpckDKUHn4AL9nHgw3Qxw7OkeHHw51a+QyC/ZRQ
gHuGQCyfzfYauPJcj1gmrclMK6Tg3UajdG7ZnWkK6CjZgJx+gHmjONP5KCePzB8y5gQsZ6a2
jYGkEozcH9Fvh9K07/hARxdFGmPwmu9BmSebjYQzMKACTLzGQAXhl7NCneKYBruIHHabQxF9
6Yz7n4XGroLrlq3a6puHEyvLLwtJ1ofuxxwaiKIrfOB0h0QVmz4qOcD72u9+FQ///I1MEzAw
XI0JD+1nR0QyqxVqgnHP3d/bBGZ4LDHQ5rx6gZx0+FyD/T1y7rdmr8Hu7yZvZ6Z2Ljnayg6Z
zMGOWsIo3T2Lm0vj3ii2etyUiQova7hzC3rcE60QeOKKSNeNXnaRmZxMKifIzf/MWw7jK9oQ
xj9OC1agPwIzWXr950eLmQGlBh7tDpYTuYXIzjQNQBydCloaFE0EfdasTQp+q3eXUaHp9xZ5
BDBK3cwjcvo9ffFuT2oJ3x2/69q6Mn8TfCQVWonHjYRqMjre4YLi2WbGJAol54A6PV+XJWgo
ZnEH1a6emQYE7S82mosG6pCniqdis8cA958rzb9TGPMBcEktFeaQd8IyS28yRNYSejpVeJV3
iRWNi/piXnZtZRx4jUyvWneJd+fJpbEcoMjIaQs6PaPupbbYm4bhFxEWK48GUwrAAXVhrFJ5
HH9ED4OS63sEWUVqFWVSmvEdxv3GNO2cQhAmAC0Oj8imKn4xh+k7ve5YBEofMFPCNub4GWD1
7bob2af+d/cXus/LyTS6yA+Xw3U/n9PnyfymVAslso3BwB30mXFvNcCNcBbar0VQXmuWnp1X
tjGIIvq7WpbRWL2CLkVg50iquR52IQZxR44I9wzgJNQomq1YUDVNci3c2mdlX2PnyyTnRG/n
PwPYKj7eEtCfUbUW1lczGHLHgCa1Ucf2Uz8nOiWra1I/9iSrKTTgVubdMCL4NStyMdcX/FoG
haasz0IkS3S0YtdxyKfejlNSufPpR/K47pug5OIwODoAjpthux4XXZKX2GyT1GBGyI2/JmAW
yFKqgxpThQSeB92oH9M90cvVegaTj0gqSkjYW38P79kzv/myJjhmJabti3iWuGqiEcXHTaim
nRk8KQaZaTBdwN9P9uhurt582dnZDycvhyK78eA9lpv2WPX+VMaXTntZ+INpR4oO7+fba+YK
/UqqbRmmo60KSqTRGxRWwBopZ3PWMpCaLsTIcIyxgBmsAf2Ik86CupEmL0TVyL0+e9eyarMm
rlaldzrbqLUUpYdizyjNEcBkLh+/wZ4AD3dybo/m+uKaJez/EeqdfaIZrHsJ24m8aFXUGEsc
D9k4lQrUg49NwVrlKHmnHNfY0YMIwbyI7Tvz+a4RN1/FlsyIqivg0tcgjddD50CGlTEyJcp6
5ojhAxubUm9EW91kY125TPDiQUZ5WexTS+bp64oWVLCdASlEGwzScLKO4pHvzOfhrio0IUtV
IXykosixSqV0etRdxwa1ndrvxEmEq2HS4GlyVI6Z8+1igMWi7sB7krpZFbIhCClzbvkbFYYf
hyF+Q8DPvLSWx80dWtuqPAhpWag9RzbSchmMRuMZSto3QYWlFu8PJ2ZlgQJ78HD1pM+DzSII
gIS8SBzSM7Qr/vmqKts+I2d9k4whpkRnrxbbeozbQwCPwc3JkecljO9wFNfmVI+yW3gICdgx
H/1xZh70bLQW9P0kXdHQbbPRl2c3GSC+xC+wyV/C7wDpWrZJYXdHBN9dgFRY+qhp3UjLG8Fe
5EM89McAI3gGRQ2ICzDdpexRJravrp+qnTdaRqSDuCA0/u+NRT/JcopwOb+lUIObPDnGJmRF
xPdjQQKUOk0rZqUMD83GmYPB68c06Yafb1z8RLiDWqSvtYToxFhSXwPlRAf7TjSDQ4/7Abw2
XC9Kpx+QpnckJtYAtaq8CJiXpzhq6UVd7FBLD22rhoQVuRmJLEYPsl1XMiA63Dk+KNg1+uq2
+0nHCG3npezDUY6/bxgHX2JMu3bg/k7hzU7Pjx6/0Zo6TgAg8sV1qxRY223TlZEhvk9yIL6t
EElP1ZBNeC4xkPYQNSEn3xLQBZb/Izep58+qQn/90Mo+SRvxgp16ywmGEJfSzSrS1heF6rly
uXTCvDX+3dzUQp6Ge1FoQFKoIuihmvnciBi/R86l4kHDnxQ4BXL7psRfv/vafvlkmc+8jEU8
Cyfum3xE/MAsg0vHrCcBkhsYf/IXRaIzAPNispW1cWv5WHpYB8N41o+fEsm7Fj0uDCp0EGZl
lglILyXOX8zkJbjiAqKjmUR2dwcL7sTQ/oBRnkjXb80v0X2QiwmaHLjrYJpSiYhYpSLCw7UQ
vEv9KYHWKFGl9i/3rd/XgJO8Q1NF5trS5xR9Q2ilLWNKPIwE3Xef/fAB4qWa7e4FJoMfJrXZ
CuhQpI3mB8XjUB5L895Y7SydAlSLwXyHrQSB6wDzBE5Xgc504I6SK18EWEYtGTfprSorBZM+
uGYDPA4nuQxDN+3WnTOq5SUJ0cFmEb6T1Ucc+Ur7d4vDLR1pNWBiG8NxxnL4w06FgMg59FCk
MDhg/jK4rVavZWC0iM6rT8DM59ju5JLvNmRp4Xg/R9qQ+4ct9SZRiqY4QRMoV1ou6MY8KwjH
5CAbgrBpdhcosF8LpnQ4HJTjwIcw/0ENTayL8UbuoN+jr7VaC8bPkKWlyycMI4qSgX5xvL30
riqbjyVuL9R3FCrwSuXBW8N2PX3RQPHH0Oe+U+EDoLUFE7YlHWGpbv+CUA+k64kn6nwfpO9+
lU31MoVSCD1LL6k2aRPpvhGo40JYfoQVjB1n17yyCcCuW0vI7wuG/pwpwfYbtLFWA3MGS+8S
fFk1vex7nJBIkkpiLg4MS/MzEu5Q90va05h1lnJlYgL7AgUYUbj8M88w9N38CUXa9WNhCMvz
lDOQvEj8mhGCKMlRlqsv0NBxb2UdvaDcyJVGT/HY5nerd82l7PJqbuSZt3ZpO2iXtGTMM8aY
zuh3DyNI5VCXuGWVDZipdVXMSw8RtSu6sH3lJcdWQrdbt5ySItYHim72lcXmW2HrXpBTI/K2
qsAGrT/yCDfFJ3CSDFY8FKlHdX23jGZuor3KR9CIHoFocWvXURiRFGJLBD1hHYIX4QSx9jjH
MrzmYtoApKsZ54J7r0yFbeNNi1POg/fdh305PfnGjApazHOZ+2TI9Oai4AorCzIkzSce81mM
SIdO/iHAbO/+/99wuxYzy41snU/C1+JlNYpBGasilIsZW+4MNzoZPyO5DMFXDoLrvQo8zDe6
hYfRxATTNBaI4xfqPwB1YzhxSjwTy7MAd99mczFXUbTj9E6za6ynmXVt3eC2JRX/E3C928kp
nrFObD1ADpQ/vJIj3Wy99k8to9tzXNmtOgw2WnbUybAWvGRF7T1mG6XwYzcuW4mnbKJL481L
IscLOApn0O7ko1EsASpgjaWI/anhxyiDyhfWV+Z9UGMGMANfuPLXF6crRl4uyk/461LBZWKl
ZtBPMZ1igHMr/8MA35QTrN4evHey8NSE24udvZoxtLMvvkgNYtKhBU6Iw3eBv2NZxED/+21Y
VqYT5RcL32PAyT9PevxeItLKaa+U5YfwwTOV7JMF+pSBPjIntilRhYJQaHQBHIA5DGqo1tdV
xUW0BbADyi8g9wKWZQP+89SZMvcC01OJRGELHPW72XMmBBY9a2TDDjX1mwWUzZYldsnQZ1qK
UAyfOoH7CKTqqcqACCW9KOKx6mkNkK+52y578JBkq/PhlHP2SvLy0AaIZEYsL6ruck3UX4op
Qizv9d3fG73+Y+VqD5XIap+8DeTFusUJffvZsj53knhGCv7XdEeI8eHwszzjenh6ZsnFATKr
gSnQ4n5dDzwovrOYxQFvTFPFR9SlH4ah09KrFFBhCCNelgs85dcFwEuVSLPt5ZTRt6FFgdn/
GNtoOeanUXliT1hVd4jlHIKlAyqYk/iZqbFk9cBzgxJp2gDKRAIbRbNj3zZQEnoFAzoSlO/j
d3UWy7nng89PCMRW1nmbIU4TL2Z/Wxjl4q9qESE7r2WW+jMAxX6znxyllfp515pHgDIpoIU0
nZChQQZfk2ZAZ4b1bUVRCy81LDEj8L5KeKvIdvVD7YMBjXjCVmxjgQdwTb8NzF1XHVMZm8G2
+H9MFT9Qv36s62YGyd5fiL3zo33qzY/p2E4koq8yQcErPvQzHly0QlVYNk7dHWy0iNCk2moi
lmFUZ9uzYTPx/3W+JwP8Aeq00P3/70MDa7/T/401qRN7azmks28gmAuv3oexSXGPCiO0HAsw
SYYwqidISRsM91phMhdDKhzxAbF8emfDkTWIXT4QOFO7j66pxLyzU6u4OV9EkJRf4YbSpd2h
HD0Q4ZndAEs2wZ9TOQf0OYpHPmdojv+H7kTrYkVRwfc+4/4jIKa7bdhjvjcN/pm4fXoO0Mc4
g/dYp1Fu3kutiAa8wwuETK0+OeP15lGuZejceZiDQ7ffEHrozFxLZs/EgMDRt+kuoKfw/G8s
i5c43OhxeFmpjKI7BlCuUul5++JFguaMqyyS9MZPy9bYmcab6XcxFjE+Q2PitD3myyz7en+5
M7k2DAhAmFz7y9FYOTbLwhcNGeZ2QDXnf+8MW2T+m9gWA0njn45f2ucGkQkmjPj2//yv16N5
XE5cTOimYvhF7h10syLmBPnjQf+Aj8jKwkEpYr3WLF0ev+1AyhLy8oMiR+WlwxRC8u2hj4vK
bpV/g/qPVa9sFMFbqTAXhFycJzQ6HwX5f8nOvt2/9yeg6f6Yth+m5uHMr6wyJIyE1aj3Iuc/
5O/jazmh7dktklAVekMSEhgXp+99Uhen0mbWa/RjhxJUpO+j5FdDum6Eeh6RIpvtgVpXaggo
Kj2gg58oR44JLuiYB2wQCLD96RlTuulcPNhmuRiq70+cX1atZJJMmOJECCm3hyDno6ePWCiv
TujgOEgdNgGhuQTb0iglyqXbdNhda6xLcNkGb7ARF4QM1eQ/omyjGg14bGu0CkN5Q8lg1ape
OXw2IHX1tMnR2tJbo8BC2f1qzK1LuZDlBGxwwVLbcZOknSRO2lrAq7wbkZWMxGSI6bQKizmc
1lTt+VA5MdsusghR3li3H48UZ9Djsuux/s2vty8QwBwgzQygwU6SB8Opi4v1282+Fhq1T7OP
6FhZzazIkusrMEKHpIxgucCn8GM+v8noj3b3XUjNkJajCpQtXvliL7A3lfEdGEO1tmKSa6zD
T03Iy9kS6nAC7TA0bVB+XyzYDIzTnd3E2cvi6CF4h6HvTzpo4zwLsx/4IK8OG2rF390JKjQ+
p+qCQ/xSLxfjDaxrJkRv5h3RcATzqJdk0jp2BZjVeH7qEiLIpax23XBagSvlXvfdei1HbXC9
AICuEjLLP+/U+liPNvr1IyfooJbVvfnPyxgqlIMzALvRr3tqTKSzOgcq8yKlwZNK6orSs28H
Dfi8WSpomtEsBxBcXXemQ0WtFwolrctgbWIYxhotf623Yh06KziODPm1znoG7wdmDZSqsame
tcc8kyX++X+d4RjjP0chtktDo/za2arQutE7gzhRfQ8YaUg/dBx8iYNPT0gG40Ilfqo8X0CW
UraEhFwcqchAuyYpI8Jv63bIwbn4g8wjZBttsK+VWt4np83dAeQz+L0sDkrasEeF6u1iSDNS
r9WGhYPTWEv/ydPTVmVCfjH73Vwf5uTpB/2BowvPPh0GtmBYdieq+e3qGV38cbSKzFcuw1sE
L+gOlbR6GN8ha9e9M5GGvlqcWskiNKktZuJDtCoViJVeihXKE+buhT65O6IBOHezfoyDMg5w
I+fg3pFwp32i9q+LGyOXi5/mZwtwTE0gfHXYgIiXTLldKhb7No8dJHTPfwG5Gpky+rhdegv7
sxdJGGyjVXGCsf3CjEO/mN5LVxC7AOmsbhnZP4Xu0KEGlrjjtKzsn8cmxRpnwQWa5plFOHWN
bZODZlM8s0xgx+CUmXuPOUbj7V37rzd/RQ4UqDxGaynie68LDpBPtwIuR9cxG7lW41IjE9iw
3swtBA07re19PYZ2SN4wo7EHCzKbgrXYBC6kM+Mca2lB/sA0OuQDUH6UQULxY902hTZfBrs3
POxu/GDBeQ7VC3ijFcbuwCgGXM9ML+RY1hd5cEhqrm+K5iqFKg/wVh6y42OO5kujgdfyoVjH
W1RHuuskCEho3R/SedLOLgIurNR/xgE7SkMTeaPZLm7tPrtvRchEwbmnvG1MnighwlEurwx+
wzwDa3NInMlwmJxLq+gtMLVv83kDyJGVLF37jsv0wJdpoylmIvrOrTpTUT0Z9tuYrYlwZSE9
rnLd7tgUP6psm+VYNE9BJXnGV6EYhnsZ1/mApN6HIgRF4GUROBWLYrdKyTtdd+DTQXsimoDL
+pHU4LELRKQxKjAcWQWZzkowl/cVPgdDvxUam2B0dQTpcrtPB7gMj7P7VhpIKzjIJ7tkQh0f
P/oS4XNC1LjEn4LbYi6MW7rB2TiQdZUI2yiY6UL8OyQQcnRPs38NFP771iMgtdy1ZBrTzkk2
MZGYaae7D4ugsjTKC0u4rhrAvOPCdAtrWdk7FxZMkmggaRAm6MtAWeMRsgH7JsAMddyx/cTW
oOfMKufOewMkZpMeip5/F+S5PlIaqEX1jz1mA9GXhNuBXQURAKFrkyGlMzTHS/B8VtC9eLad
vlpT0oOIuMcn7R1hNiZ4w8ExZrgUG+aWBhVfKikg5jm1SRVkiMoj1Y7HZrZb2gHhGtF2pB5+
jrJ2mER/V6uqX4NnxA+jXCkhsvjrZjjby1PJnkYeRIPZIQPOh7kJM6nUoMlYUscvoCdvHaKJ
hbckfioka3EnCcHdjmq102KgQHVZuaPNunSxJu973CbAAqzydrqpPQjyQaruf3juwGjz+iek
LmF/U52kzQyCrF8C9qo6fR0PSX2CPLhdbB2l40sLr7Q6+BsNZY6WQC506bg/8DZ4N/Br1J/6
55TGp/D+FInkkQjZ442m9RPhu++dVUmD4jIUVriAKV7eXxyRbbk2dKafg7uRrTZugwvPkcd8
sZEKydPa9OVG9za9PslvtG7INNSK1IMeWzCnbOYQuqcKgkLjodl+NrOmfTiGiKSSX/fJdzHd
yhjeIFDNTcYoIabaknhlIIO10rQQKplgYSMtvFFlWUtt0ElhiARZdedI7762K6bBX4dLkh03
h8Em6w122NrymSrD76d69MwF+JYYoh/2A32Q9spt+q0tuz3aTgScBNccVcbDLV6e5jBL2+AV
E+ac+gi3gflM90ZOjbXiyL8TivYkVYHPLl+vUpYTHaf2VSrKIxdrlAF+5GXjzwjaWHtE0Fng
bYsfEpdqccvwehYrVwRyqQt44hr5nWiay7c8xYWbsO39RRc/IbIrrJTOaCh83zQMjVZnrY1H
f5Y0zVmezYGydECnmwSBZ4w7iTWazT+WydlhJoNRsL/wrJYSqk/+HhQrcVus1UZps3Xv7RNt
QGOxJGsz9Odtm7PIEaymEmHWVNbRKfUCIqD+FFpaxUMgJ9xJrglTDNRRV9fmUn4VDaVQ9NCL
/RtfxINBw6mRGbUflDC7RMVRQP0zqnmrMNtE/DfRGt6iub686DMJuxurM/FYWXadrbYhXVa4
MB1QTzYeq+YMrZha4C+olZJRa1xPEqbswbwdWz6C2yXig5GTAsLFsgE8cGj4dG9r1KaJmpHY
5d+vGgQc5/OvVGOCjCWF++0//Qwago6iNuoH7pbixtvO/EwnnzSY4+K8hRKJBEYvS9SltDYm
aiCFGHjuEfOiNaYIyiEdN8muhHFvwXlf8SNMCrs1IfAiHQED6LNNGDXrlrvLrkmUF97u5uo0
gvZL45A2T2DVgem9y+2c5P/C75219mZlRYrKAmTOgaHRQrqYjJk79qe4o7U1wUcaN67VmnCH
MmtmTUkAATgfkHEnXAY5TopAF8XgpBE+wxWb01G+Rf/kecebaFY3T4nqsjMuoNStDiDlZ6+R
2zOSDp7FAOZiskZxOAvgsfBll4IZ0mAHFV4pJbMmHHqFZnTxFiNNOHPmgH38ua1Y7ncPz9vN
6uVaY3qmM4afPlmN/oE+JYjI+cOK614GyQO9lPG/+4vfm6d4NNd2yazvMNtGDBeHWeEI6p9k
HDpiHWFoq8zaVfGvMN5sGy95WAsikwaeFPx0BGhIvQ/Au8huRsi7JANK5s0EO1/4H85FYUJ1
ZXNOInbkOFYj6rj0zZyAmHXzI56M92/JroU1eEOoDVHNmbQYxVsmfWLRgXtrX7QGpZyf0ZF2
i5vIrmrFgf6wpyE2taajn9R02/TL9DvoonAw2atxiXHW44T+WYgFq03X1Wfr+tStsQUSvVup
QWNwyGagy7z7AtWFSI62I+dJbV76uZ3ugCsqwK/M+0m/58a0MPPKZhcTMOolEK0O4u6hD4e2
H9GFKt447wr4Gbj1lWO5fQVcU+rOU3UI+yURYF5k/zmYuJii1JMwfKrD/G8TtjmLUaJ2SBBl
Mh/MDAryfWZ3NzQ6IYB2/DO1mwfrZI75lyo3rxK5oOrhJ1jQTcxpGdti46c3hHTG3dZQ/Ige
WfBecgUCFk7L3s/XBT34eUrjgsov27FlEXBtAjMMWW1umijlMNBsZoWUChPyZGTf0YZF9jNB
ivMhjf+i3BxuYaok3JOYsND9E2PyZkOv1yk1XPWGIQ66NBzSP+ipT4Si1jmU031r+w+HGKJn
x4KYIo0BMNYQo4/ZtHRBahp+JhpdyaIsXybFZAth2xLVRlZugQhL6qVegvpdCAk59wH4n44v
cHctsKoHs2wfNPqf0mHRGNGCtJQu8J9dLXZXK8S27NKWZxt06Gm8l9UkgMoWlwrBIpl0b3A+
rnsR/vjRrrUsolKaVdJg078tHYbFSXokug3C1x9JVOOzSZUHBsUfCJrtasWZxx8PWwZwnfor
jTj7OajoI9r+u+h9EyzBwXmSZATaKSeYTvo5ZRhVOQ8MbnMtzRdfIVjzC2x/tuxgwj3SQjzF
CgtFifp0NhmitVHerbI7qySpVX62hbu6Ptw1kTp2k9Bv+mhXfvAQtyLKJJmcM8+nzP3hPtbz
y2J9T6nx/wclAkDQq7Hw3/rT618wY7K4J5wsz+cbGqUIzBalSIQdVKa2MeaB+J4X45/0GbTU
aDSRyygg4ozTuEN4t1n9EyIpZf2Q0+d8TEJ9qh8xEz16nv/VfTiNkIkFyOfLdZ+HelRzUWoC
bk/UbjycSq1DQaja9XUzh1O6OL8B1kLJtcrDlQmNZRDeYwNgtiea5hNtv6hw1METjW/eoENf
3mQAWZcRJX5JzAlVsxBfxqmR+HXYL5kap+tPVcBgAxll2G4caM0l5rjDj7SFKam0wLN+kZbj
FMUKkNNvxpu72dnJ5soxrZj4aUj5CyPtythF/rUjwGLwLzMcj7cdIZzMzOt5RVQcJktb96lT
DPa4VH3kkP5zvSAxE4C+HWUk+eJY4DbbijaTFud7J20loywD38aBg9caGOoQunYVR9zk2h1h
KOTXxianWjcKEhOvwtJLUMQKRfSQYqR6JX5X9ExpncBwBpj/h0f1kkZ3xe/y4xvJfoUFN8R0
IDLo6NdUl4e3mgTt7LG48HUVCYkpXXGIK9qZTyNwd4ld6YhxUO4cpaplKT2eouKCD1wKixvn
/09R0K65t15aFlaXtdMWAQi+Mjjl70040WEjuvp3glXfKKOm/D6txbmlMnLUVQ9fkHXoadKc
5sFrs658Pn4fd4y2MM+wH1shpFkN1dk/8++TsZArHTtwAEmfK22XFcKKqDK6UryU7Ka/Xzg+
9yzrD/mqIM20USqrs1x2OKdEFbkYmW5eogU2QiAXF/TL/7tSJUUS2LjTP0mzx61KFn1LmJ1P
yQk+80FnPja3EXF6/PgMzz0d5SznTvAFBBhJnIPRDiHALPeDLs8AuSys+Qq9re9J3syRbk57
QY1y89dHdXn+PAWG2DIHrDKcTZBCM6wQ1oQ58+mBRQf3AVbCIUvpdhMt+iNRMiLkEhPekz2g
UCVUph73caf4MNwLsF1uanSsSXUmIrzNlNojPL624fEiU+9K7oNHpstIRqA1oLju8UunkEE1
wAcx2HsKZ4klw2VhdLkFD1Fx9ER8TrTFEpwa06RllNMnKhs6Lf2NVtEPuKBCbe1eYLAkHdeI
Id4CIsG1wLWj2N4ZEkEbG+GuK/1F0FeONYN1vFC8EaGCz+Hgdi4g8zXjvrEfNF8LqtYRqWwF
Rarm0e7kbJZxMkXtCSF9H1IeUku1YhURqkWTiPbnwXJOfBU0Gw5Paim/OtwugVexarq7+J14
6TjSh8oWWaBgnhN3c/z4MgqpsYPinbpJhSJZ6KWkXWrsQp55p1JamQNH7VYe1otktn0ifAag
Y9Zia3IKHMtnQUMvsVsH0ak7M+utCZt7YDnzgaeRz46Cey7Be7nThLLsaLZ/JXtM/YWcaAMM
bKd54P9xoWdnpRgZptfJYHG5kcbvi/fK5m8CaoQ2yrfUoy+NAwgKFC5bIIB47NkRbr21MxsN
ZTcnv7ZQe13BaWuOAFW8Au/ZZ6mrkZyl+WQfr8pU/03cIjzNQ49i4IJUKJOSObSYPLFnco5t
igMMObMCVhAj0TBB4H+IV4YAAZ3bW0YeXHWSsHweVn248fmZO608tLBnXr3Fw7Qg3iOVwcOK
yDqoQwRio/T7vjIjD1RbwmCMcW6qwTmsHoSK09pZggNThNZdcZfLgKF7X6S3I1xm6j0kO9RK
fb9307KmIvmphaK7zjzi6a7g5woZcmvHRllAfP/wvqKA4P8nNrM4/HAdc0qBp+B1TlSn6PlS
XAer1bOsfpYVSE3jKxsHJXQzLAb9bJxptxP37O18RUDKDBhIvZ71YE9OvFlH3RAx5C/gjoj7
OPjcXojmSV3n7uTcOgm4F1qsYmnpW5ycxRawX0ucwz8gLWrbYuoGh9mF8XcdOdFFZekD6AZ6
Y49HbI4RWg0L+kIdkp3AF5vW8Ri8MQr6aeGeB8l3tdw0wJC2dxz+no+aZgq4mvK6s7sYIFTO
Y1lbKUtMazc1aVDzxrWuZd2nTddJB2uqhnlq7nIKGyt/EY7RxZ1RsrnrEFbdHy6ZFYjwiouu
sq+f2gEyR/pqhM+QoCeAEdOPqocWHj+KHl84fsccGvX5dE/uY0haM8ke3qKSYC54470e8lfj
jsR8SBmX30TKD1gxCLH/2SIr72k8HqpshdjPxKeeg5PuTINuZeK7sSWpxsIHLm+2vQ3sKFL2
LFsDqLRt2BHnZ7kjMbZFwNsuBbdFblnSsmsuqwAu9AzUm9P8aDYZ5jzd3I3aWvLMyWrsmG8M
lvH9/y/22Su3k0IQGvyFqNPShLlpeZ/kmpHBb6rHTt8QR954+OvZhL9vbeayqanftY8daTTx
hHDFK9utvVZWvd3MZhpUm6b1Hb0WpPxsw3H82/prDAtXlne+Eh8l/K7pxXKkIbIZ0jBWCyks
+hFRB737RIjCx/y7eUNAN/U6LqYH5Dv1HAo7NIlGab70xv/dkIJPiKd7SryUwFL6rcJNdLg/
r2mQ/HhZXGCUkVLX1EHx6YzoqHA214zkV7iLX9g8YuLc17Um48LBh1wKGMUSGnj9hk3UkXup
dzyhE+h7Fn6i3dAO0pwiu+OIJtSqd003crP3EtgPT42UTnx+R9WYxgQ5/IjcGS2LVTGa7byw
mKgQNn3IWosT2kcSAP83+yOgI2u6eOMx5P1jQkhIkN2DL+yGy7pgQVnR2fPxzJ2Wv8/oMP9r
f6//7itH+D0WHrPihQXkLfOZqOh4zRn7+pHZBq3IvPmyyqCO4lKx5duk7pktxuL//kBNvQ7j
5G4+d/EtWkznYpDwz7fmbm08DYuhlJtnlVhfSsC2xThzDPMatBqGkZW/P/IXDf1c/ByOSbtg
WoLVupnrZnT8uSI3Q0By37BPY+2rBnzC4xuOIyVYw0VU7e7m7C6vWtXvrONW0BC2IiN2Vmmj
jiJc8xHlzeGA5puI1WFIzsfnW2wN29ru/fpEyuLH9aC6k3vHgZDBHsj+zXQnQ2tK/WqyvS3P
xajSXbxig1bHy7AxJtppb7ICkADQKF/iPg9jCh1FOkRsvRTFkuPS/IncNATFZn4xJh9pu+bC
5mdNWV70BeSodYWkuzN3oCxRVhw/csb+2mMW2IxQE3o2IjiMS7VxgT/3fPEJnL+d2ftU7ByK
RXluVFMxIa/aqi3tw3b27lHYvzZSUcCr+2+u8kevv18Txzoih7ihtJKwXhJ+JXv8G0lM5d9b
4Fm7n9LBNOzdHbiqLvHGWlhQUjq/IRKyjVQbxlIwP9c33bjgfUb+MHZb1ao9YtsTArMOGHif
zwKpMraGA7nC/sY/pk/6BYG9oM91fPCjUK/pS1wJMVtf5ExOKmw47/s00znBRZLSR9LP8jkP
cp827rZLOqEL+vFUbIg9oKFJaY32aPq9wP/DIh3/pSWXGQZfNopKJ0uonROfaxUE8TmGqFWx
el+9MwhoDtlvLm+FBaClMiVo2wJ0HDVtF1jbR1vY+oNxcc26TVcSN/4B+62vxR/yS7g/pWK4
k7gyrq+g9RYKUnjCP3WV8ErOiNeBwfhlWMxgqWRXLynnTQMUD9Z1yc8FX930p58mqTOLs52N
IHSRW7Q5EkUg+ffCba1KWqYvQJOMbXCGuP0YxOs+JdZp2p1RfXyazjAZ8SlXXZ3EmVQZyFmn
QsF+ecwwF850yuRGO2O5Q5mBbcmNk7Glrl/GuDA1k46uMn/Rz+7OBJQ/++3ceIAUgMvXrLFv
Q+hLbcJWj/All/aHmh11Pci73aqyrBzmbsPtOjriJKjiucTuyxRc1aDO3H8ZvAXJeVlxBTc5
C2cuPAav/0l1SZ39LUW4GwJQiP+p0sGQY3FUjFoOEhHORun+/kvjs7kEh0/2EQLABX3vXzVC
PUY7861h2iw8bNP4QNbclt4jIGZkzR3WxN1w7J27tOJVz3MuabHlsFQN7mECUJc3tcg/7P/C
fNgkYtEndxPHC8nhpjMnny7OBTDg4m8kE1UP9KUrWQZcNoKZRRKPrPRL2B90VU99XIun7Cjv
p+g0xDHmpNZUY0TmiB7ssx0S/Se/MuWnxP6XFC5jdMl+88tyoqZXsYp7GdcEBxFRYjFTZY3k
QeUM/K72mmLmgb5knfYnUBNjV9rWC+BXRtRXThHBG+Dgwxns6oKQkmofznyYUnuEAz9643WH
CgRabq/l0cCgc8ARK99+vHAMjZPHTAD8s1dWYI89ASYrFg1+VPMMbG8g/QMI65BJxUwinmHe
S76E2x9LzsaECIPnndvzdTe1w5eOMw2UEhFt0GRm0eJ531QbZ4trvAIKqRv8P6WVeWNy0Ms5
7wykRV+72rg8vFysbU6FiHI4tCeolo/kssGxF3SXNuHK4rR3q/v5kH5OSLM0Kf1b5wE780OT
M5FwbGOsJ5a8y6StOLW19/OT2WZmjxTFC9aFwgvEVipGiNWSKqfkJlTqWsfcd5M0URe6jIXz
WCfbPreCOezVUUYdFp0/QVzagtEvfQ1dcGKinJNJ/CWpa5NJoZpB4zAcGIDcfzFDlY1zE7vT
mpZ/EJud7YOXnp2ONhqCU9K4Ymi86/SrN7bEj1GHEYQ2BMHYHIKBR5vlll38KSZfLx/DHCkT
S3CIZou+wGZkyi0FfStij2oaIjCYxWkAzFvTkfi/4x80X9OHH2vtODvPSx+oLjQmYUlHKUgI
VregR+evYuUWIvN5Vs0pYu/UrCKPcQSKV5LaMZCN3djVaXjmNU2ApHnq4GYzRbT2jYzRyG5Z
lYEabo4ETLxp6yCSJnJyFZuTl99r5NwMhNC233IyT7+ExSKjw1Q3Q4rpxmUilNpPfQHIp9Si
eGl45wWrxXXh6ojFXwqJF9moAzIe1dd4UFiRl5bENLqVUKQA6WgtUkxSrIBV+b4hcwH8QgZb
t3nYY8yqaE5shMqmqfO961jvqdV8O6c82Ht/KUf6xUXcYSvAg2jP2yrigoWdxazCiS42IxNO
InrDir/Hl24IE6ZS3LzkdTXi9gv2GKpTLEqqmoTs8HI9/pWIKS3kvaZB2ozZ3spwWbZL8zm/
/1Grrhhkd9UC73rZlls0MO7AgXlM1J16V0MA2pPLJ38qO7tvr+bxb1Be8VxN2oLTdqeHaL3j
lfZ0N/3cfJkIlIcmwkKbD8ipKjR9RvzPNfobB/0SXpxTMpot8kSn2YH7rLRv8kfC0DGK7g6n
NBAuAlQ6wXM4UoEUZn64GFSGgX8fy9AXPvrixeVPJ7qsPVGxt6kFR1U94kexuOK6VUnytU0+
yYLepkeWAOIY/GcDT9wtnAdTaRYCqKoDevX03qzdmk/DB5bVeITGFZifsya8ZXnOLcbdTOXj
olP7eax3rE+XJx+oJ4LEAke1JTxXWg8Yo3OumDYbdDszM9twYaaEbXvvcf17ui5BzsWHJRGk
sD+tFiA0/Z468clK89ux1yckfMLXv8icIiRRI2HqEsis8zwF8fvxhQGi98/XZ97WUfUrxcMP
2uhWzJSbobW4INKZ8mgPL5WCC9PKkf5tYcXK/ftayZ8cK7Tx+j2+BeC6TBc3Q1xDi2MvlI6C
wCZvKu1FPxBA+0j4ECUvK36QxRnbl59ysgGyKmFgaNIMt/hQv524EpmvS6Wi/pHZNE0Gp9gV
id2SNwE0/3F9NnGBuXHztyu6xT1zzPPwT8g7jCpktpcpMbOhUXMR6FxjvgC9GdFs5ZMQkKqU
f/JkBIIUTatVteIv4slQPh5gEtSzBTQrgF/ILp67+OU3mG3Gp4qLuBTppDnUOif1TIvA0Q6d
zLHzyww3J2ZzbJZWzDruiDwCprzj2j0RxhBri0YBY9aBuwonF71FtzpkK8GxFyEz3L55bAkG
KcGtw+rjgTwUvLne/SDBjVS/tT/ZKbKH7L2EqxaJaN2y9NgLVmR6dJsEWDpJposPQht6cmwv
ASya8p1Sl86BCpbaqAeRieI62MhJoMhhRZb37SJlS5gN1TD7If59sPz/ZN5q1XVsS2YEJr/m
W1K+QTi8YU4K+qKmY678wRpBj/H4XDdTC70ON9NZcFC9mu2gadQumt8OAalwbQ9hEtyavgC0
9HN60uMTpCtJT77/6SChoOc0WKJHzkObmeUb+laLABqbDKkCXB6MlW+VbjFR+TKeYoG+yGwX
ui126hkLA/4QH6/Z6CGbnCDOFF5m+GZ1aWzvaqUC0pvE2xCndCOjKbM5QvpUrZ6O3XfVJ2Dp
3zAk7PGhUeq7OS+sA9IaGOJ5XutsimtSLnvh8NFX+UR2Saj5M0L3/XiUwXIsvNpCbukeS+Gs
HmX4LY70hXzfY++iW8g6CfUq1z9o2uZf1S6ZU4cQimiKHas5S/KsX8adhF7v795Tg9KJnzM1
BGT+x4f4wyX7vpwsiYQvAbs056NbdDetdJLGPAeFNMK71Dio1m9DPGp7LwZtqvt72IGvkSaH
tHxQydoMi9EnWfXBBXcKgT3E5k2y+UqPWOizUAjBzceN/JzwapKvbxdGiHJ5Tvnl9uhFFy4e
DXIevqVmzlY3pqC5HB7iWtbPyreZSLWOmFoyv0H8V8KmWdksHAJ7kLoD2CEFeYU1EFYBSrzl
bxfd44ktc1zgUI4Pe8OMjjW5BnjXHoMqb7oCY37V/b705Ko3onq7XBPK5nDOsMWKb/G/6IZa
Z4eOpmQA7y8/rPa6dtpKIHD2L3a3lJNXni3rvduW8pJaUIAuxtG/RDOVlfng6FQYons55EyL
C4iHZAsqILmktdStqKk8eTAZvLtIk1onWOmodFMxwH4ALiVOJG+Y1e98YJ1WKbuflO3hIZZE
8PLGx4B10L0ZHMHYMQlC1FakpGk2Mwr2cuu7lJ0Z4j0stpfbW4H8JwV5Wy660ZwUMtJHNG8z
LyXJYSDxt+iLyZ5cArvzPx+9g8mJ2i6MvjGxH6G/+fhHT5sMJhR3dn0ovl/pa/lf9ctke41r
rQW3V8O+wvU1MfthWlqvnyuegmB2DSfWbJ7kIZ7Sk6nC4gpB/NBn2dINUjqdYPO73k9uGsa0
BfFI/U5RI7nTsasrErJyF14Lba0/z1PIV06tgdcAQBo4DHleURNkpK5xAbkvaJJpip9mif2z
qQIHWmJQGXMSDkcQNJ8eMQ86zENCVUp+P/UD+UWZaJATMnD0E/nogPfP4gP9J8/chFxNqdAQ
hTce/HB8LkNq4kefu6ZUkjXMjMZRanndVWTd4EwWL3Uv2OB71e9PV7Hz9fnvY64PGUCCloFf
5jOP/8hj2VYbB9t3Mvvnvh6sdAlHkXRKHaPiu6lL0WkI5AhcgjhlYhcwxSz3h5fGt5vq2YU/
CqWk57lL6R0yQ94sh3RqCiYhZZhmwL8WRNiLdV03LTxaXliSCcCuGfUST2zUVsrl1jlC/rSS
zm5jBGDfKkhorM/tqftyTWFUtO+lYV9A0DhhCvUP6kB8o3WHkyJ4PMf6b5DXmFuErh4UMve2
t/sfUjJg2+CrVBSqiqtrGd/b2IXJOczewA/BrlmqUyWy/Gjpryk/s06xPwPJzIG2WC8NnOzx
FzLYQdtKlF8A6xeLZIOEy9rxPB8nD3vcURq7qbkXkvdPDyWaHreUjX5KMOS3ixUAX4oraEOF
c2dxIFGyel9gUg8EPbVaDmoiaveoIbJWs4V5iD/p05l0mpgfWVvumMPnBH+zw3eLQYh03LcQ
c5gjVOlptLyBGaDYZ7LWbIEVsu+AgV5B/Gkcb4kPpuEg4lPXEI/2PtURbBxw0bC6rPC0hAU4
vE1tzzPl+B7JU1Qq7hiLKp/kZV+rm5+D9MEdkZS/2EuuXKoc2dEO8Z5U7oS8vEDrFVh/iM62
9yLYqVBOWQyhbNaZlcosN0v0vY530zE1bXaH4TXD5/sBn3vvyh1Sb/bNL274GpQLXt7gCADi
eBZpPJVOGfGPJo/jlK9ZBNW4zE8q9ASilXnloId/xNYcr4FCIRsySNJ6icfk4F5rGp56om7/
sJ49Zr+j9sonrBmfSMfCEzCgrYyW5dZqF02Fb0KCI+hvK9D+EHdk+pkPf6iuvDevMPgXp2Hw
fVs7CtTbSr8pHBYgQyM6sfdcazL0ef8xCJY0IXta9j/6Xf6N+r/tPJ6ivHEFzMXx4+Kf0wPW
8L2VqXfZTL7CqcxT2VqUtq6xibvplFbl/oPIHiNvSN1hasHsbrAstXXkKmpZI/u/YF5efFJu
QlGXG7wxaolAZ0B8XwlRWjXziHsluRU6c2qPxlaveVxFrvC///LPO8sRJIuVazB3bRmbQ7TK
5QoAxCNuTFj4KXAAkT6F5/LEKPKJ0+z7f3CIClt9MKkRMsnTWNph+wEsyNa18x8g5jIXLZqy
rJMxcXbp08atINBqJjkq6Mefc61o21/gj+B3tqsOZH5VqVZk2TnWZ0+GnE+efBjXGIqURM/d
PIV5FPx8obs/aJ9rQszUKJJeIOuk73GOFgXD5Xf5/geQ4OMqCryaTUWw607u7gSVU+2lNEFp
sRO2I6jwjRyE9ad2dGBzdIeeEBSyEPKMXjogJmLkpP0hD+T+yx6AAobfxLxJbA659FHzK2B6
sfdEFd73+Vj7A53oYQvAYMCFI3YIiFqrqcGhDQzOoNQtDJf+Zvz4+hYSEdaP5nI2o9Hkqe8G
sAW8pR5tCHx9U/rzGQS53kXGe41jHQgcxOPhMzt7u7eHHm74Cohg0YhOFFa0zsZKNXyTK74+
W8NX15qAxx2rKt7jRKM4f29cJXpRUWFt/OxNeGF6jFJJHx/n4oAXX5yKgcRQAQI45eKoKTaj
RPf4RSJ1jpXgt9E0f6ahYXqMRpw8iGeCHqfs5QIyJMf6+tPfTKDKXQbPsJL5FRXOzmXsGRwg
rinKkgpXunB1R6pYnr3gPtqn/YDWBkGzy7Z4AYTsmSsv3g4rL9UA19KnPVV5oqWBZx5qSZ63
vuqgTqmllCFZ0Gj0hRDY6TACK1KPvlnW52ck3LWegef9D80UNQHuVVAnj7hv5xJyagT0fmze
rvxUP03b1jY5S56jZcu8hfCAzqv1Bs/VlW2Q58NLCm5W/YVV8JkOI54DCrStv5AMFWybGGZF
aDNvRIZSx6PzHknOgVFwWqo4JnnzmzqK5xWwjcAAWz5cSAcSLIvgMg6NcOBG7xDaY4N7ce7y
jGKfh5E57nNk6V0wG4QhTVYW/6IyRqKhfb7CIiMUYSnvdIiCKfMziQzkXkXN/7fKcNMpFWpg
47Hf66q4poxKmx+OWm3zlpFj5dVaDI9sLewM6CkpujQLdUUru0NYfuW34BThvb8RiBF879Gm
12kLsfKi4G0cYzj6hkQCZ+DclwRxnfeXt7ZJXxHfN+BRrKVmckDq9p7DDX013RJxgue+wkx4
du54b6qCZ9cDDl+UfLt8MO7q61NaVnWDCVNxFZ4dIarsYYmC75fmZwiw6SBVrBgCoZmXMrL/
CxF1hkPMnGg8+p8MqqgyUuYYRIS4Q8fW593bnLCitRsk0S7gP16giIxPyKNgp2uxmMbajOWq
AridQHW+ROZ2A81ePXZCn3ArbR3TdU5og+CP35s/yn7WgliLT8N+oTnzdQgHUlFum6MaNKTR
nC52IFfmK4LqlAnlD65DdrHM7jsXUTN8MmJa+xf+axOldUNLUWuYXJU0GCOC6hYmi/TZIrBn
7dlYogja7NwpxrS8VDs0nxkNum/88H/aNZz4lF/mfcTKy2C8pMlG8dZM3/YAt7tWHFoPphJy
VByYXHQemNp7oec4pPqqV1Qrcn02+HGt0OqLjbiEBF3oltASHX8x0vLHs4bhgI6vM2pjQfxJ
hT2eGpJv4RDAjetjCPcHGlF3qFSCcHvYt9klK0cYjubUntXly9SQhr0YgbG/NJJuvGMH63+f
dodUFlMR/JyWMCoP/bgHh/oPgA1DTfGKyL+/bgdVUo9xGUhB9aQNePcn1RVlNZgI7dPyOTBR
TpCwt+D+GYQjWn05R37eJVVQMX4/hseQNjBP51jx7aP5zkWGPpe8i6zmv27DzmOzCSSWF6rr
zJZDpk2+1P6tJThQD4C/FgxpUPnw0r9fuiKS8lCux20HOhXFTF5WbDnae4+x3NCwRO/dCEcs
wWmMiPMgEZbEsxEOZh1sQWkqzORwhEAsKgjKi2AJ2uq2mnR+JtzolRKqdx6tUjvaawA93PAp
fXdomPSjYqDsJDrem7YmT1aKxah1J4eAnkoBWfZy044FZkg+P6RhL9Dqlgf4Q84u/JPjOQx/
238nlcEszLXca4SxJ0w=
`protect end_protected

end Behavioral;
