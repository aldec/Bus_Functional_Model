
`timescale 1ns/1ps

module Ax_Axi4MasterBFMcore
#(
parameter DATA_BUS_WIDTH = 32,
parameter ADDRESS_WIDTH=32,
parameter ID_WIDTH=4,
parameter AWUSER_BUS_WIDTH=1,
parameter ARUSER_BUS_WIDTH=1,
parameter RUSER_BUS_WIDTH=1,
parameter WUSER_BUS_WIDTH=1,
parameter BUSER_BUS_WIDTH=1,
parameter MAX_BURST_SIZE = (((4*1024*8)/DATA_BUS_WIDTH)>256) ? 256 : ((4*1024*8)/DATA_BUS_WIDTH)
)
(
input                             ACLK,
input                             ARESETn,
output reg [ID_WIDTH-1:0]         AWID,
output reg [ADDRESS_WIDTH-1:0]    AWADDR,
output reg [3:0]                  AWREGION,
output reg [7:0]                  AWLEN,
output reg [2:0]                  AWSIZE,
output reg [1:0]                  AWBURST,
output reg                        AWLOCK,
output reg [3:0]                  AWCACHE,
output reg [2:0]                  AWPROT,
output reg [3:0]                  AWQOS,
output reg [AWUSER_BUS_WIDTH-1:0] AWUSER,
output reg                        AWVALID,
input                             AWREADY,
output reg [DATA_BUS_WIDTH-1:0]   WDATA,
output reg [DATA_BUS_WIDTH/8-1:0] WSTRB,
output reg                        WLAST,
output reg [WUSER_BUS_WIDTH-1:0]  WUSER,
output reg                        WVALID,
input                             WREADY,
input  [ID_WIDTH-1:0]             BID,
input  [1:0]                      BRESP,
input  [BUSER_BUS_WIDTH-1:0]      BUSER,
input                             BVALID,
output reg                        BREADY,
output reg [ID_WIDTH-1:0]         ARID,
output reg [ADDRESS_WIDTH-1:0]    ARADDR,
output reg [3:0]                  ARREGION,
output reg [7:0]                  ARLEN,
output reg [2:0]                  ARSIZE,
output reg [1:0]                  ARBURST,
output reg                        ARLOCK,
output reg [3:0]                  ARCACHE,
output reg [2:0]                  ARPROT,
output reg [3:0]                  ARQOS,
output reg [ARUSER_BUS_WIDTH-1:0] ARUSER,
output reg                        ARVALID,
input                             ARREADY,
input [ID_WIDTH-1:0]              RID,
input [DATA_BUS_WIDTH-1:0]        RDATA,
input [1:0]                       RRESP,
input [RUSER_BUS_WIDTH-1:0]       RUSER,
input                             RLAST,
input                             RVALID,
output reg                        RREADY
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="unknown"
`pragma protect encrypt_agent="hes_protect"
`pragma protect encrypt_agent_info="Aldec encryption tool"
`pragma protect key_keyowner="Aldec", key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
JC857JaOqnCNmsDeWCBZWWlRNwvEiBbIKtOAKcqKyQOiOFTDkW433E648nhnM2lPoVVtWAjb
t78cDdd7sEuMeS78vOSHl/BBOOJ25nbEKlokxtvEePwgaQqOSzb5yCtO6NEmDZi1ftzPGNGw
Wr8FV39q5tyTSKcW5jFtCklq+xL0fLmP5B+89SGnmsmxMgnzUbPJdvvXXFz0BYAwp5jv7+oz
gDoT9g4OuFCvcRGV1VYQsJkCML5cgJPIJb/PU3htTWAX2sW6M2x4aQlVru5WTAnvhKWXHpnC
ZPGWGrl5fBMX8VuX9LFNrhPaobU0itgaoVoR+lTp+WqqxKj8Zamm5w==
`pragma protect key_keyowner="HES", key_keyname="HES"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
kSVVfUiPt5kCFkcLWnr3usCKUXr+WqP9YuLQ6Ul8eMwuiygiQPhmK6slvjYLrJDvT049zQRm
0Y7127XMp4rUamxHuoOWrRIPbYsFkOmABdlzGVPHX2wfr3Uj/tZp18R6wBcTgcbYnrGhnyMS
g4Y/tCgMDI/57ApfVNyVpjUIqxs47DzF74e4nHw1JJp44zYnIQlsobMaN/v+NjaJHWZnC4HD
/AKo/pmXQ22xx0ep0aycDUSABIX2vkv+52hRN0lRx3cnCVbuKxO7syJe6gwKu9QpSr/YaCl1
ktkpyHYkrlszXzYa0FReLEG9I+l50wJJfx3roK2vTt6QyPI3AarXBQ==
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
JeiS+ZtA14717Sxl4z/GSY811F8MT2QC9sWwc0J4AwEQRQOJdsSnXRjoBDjKdinBSEL/y+Ea
aWJQY63FQLcNs92XLVrM4Pw8+FwgtJUHHt75z2YhJK86+ewpHMFmOel2jHmcxVVYnx/QofrB
3sJvAfiOX3+B1JhNyPJEZ6qbXAneKbDqBn3wDq6sgKrAV82E+GZXSJycDf9DqD1PwmiIknSj
UDX92vd5cHvbO+MNULEuW3kM99wV4Gj6MGbFMRpsnvQMd/3RPoZrVpHXTeGBeNQf6MXWegE+
ROrpPSVtbSw9ynT3yty5Lf/fUxVr7LipDNxWBe+nGgFfS15xgUhvlw==
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=128)
`pragma protect key_block
IruQY2RIQowTmJ60jtLfGjOCRAWR2AA1BZI5d3o9P0bPWEirkGa300r+QLy+lRn7zJhowGth
eB/jpof3aEiT1dliWv/FpGGSzSf6JQWqQqLX2pBeskpZI0o+oaleH4Hqg6cJuvOwgBPHUF0d
y8PMRH3gEZ7gxuNIJLRnxnFcADQ=
`pragma protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=960)
`pragma protect key_block
erHQCkp7ljzXVO2LOWtEm5ioimnOdCWIJqemIKrTarwAYR3mNYkNHkJikERzJDaHBlvvOeOL
2tMY4y4qCeI+4YIlB1o3qcoN/7ezG9scwNJ8V77W5IvddM5o5wRcvNSbWraSgB6hCNJQ6jkm
ESWd1dEJh6I9RubbBk3wmoZirNrliEkzE+yiCaSl12bQPW3LjwiLbA7Y0MzIVikswapx0YwQ
O2UfHDoQbbxDIS50reOM/yvyIa3/aZRBk8+8KOreSiE3gOvAQ7qF3/F62vNz2t/9qWr7gIEb
CK9x+P2/ZP89DvQIdyP/JgCpvoZPQ3lxKF5aq3iiJf8SbZNtqUkvR5K57Is3QcTsJPg30N+j
2fPIPIwS9435zZS7OqSzxH6pPNXp28M9UGGxi5L2ZnvM176jp1edNEImqfxbC/YPR7HI9d9E
TgHCAhONsBaklOW95445HKUFRUFjhw2yGosornjDqY5ENVp9GBt9OSKLirIS2ObgiESeBPvL
V9/NqYRIZ6k7llOUf9c/EsgJuh82s5nURPAs6NnyJxWgJ7+1wfg8j8h05T2uH8hI2neeSk/4
cTX6hHm092RHGKU06MgS2XFsq5QhB8r/eTcvyRwc/Yy4kEIlK6hwlS94V5cAZzvEJYd2ukvG
/A7O4kVUK+oARUkEfwJdDTSVqSSKCje0RI+9rXgWStHyr0BIt5dLcJ+tPxiS46sGtCUCc+bH
wfjY9WyZy+CPbMGIgy6NGoaZSOJgdewuLvFNQ+yydz/r4fwRQeqf/iU03RMUo1SpANijUM5j
fMqK+D6LUqK2vltUfV0dh5GdQw3eI4A145qTIi8oXfJ+prrhJjN6aW3iVJKjWz0KxZ2pj7ec
NiDfmzVcukC0wvEQKVPotXvPau6tkLefj4FKs8HvZLtZbGS2gfojKUlgqnsC6cGwdaHdVGnQ
b6TA/ThowtkUljrgyU7wQ8z/kAvveKS9GO1ZgKfUjnxlaBzOLcrdy70qSxjZNMRQhy1VZDe4
x/1nHV46SjGig5R2+hWv2bHMQqvn48O5lZkQv3RkKMTp2Y31PXOK0XJt2+osDelHhbdj9f6O
O7qaIeoyCGTTddR1UonBFyvcw4QR90HPDN3HL5hJvgFpzv0RDQvZw3iIag6F4oCb4ZCTkXpr
Mu9riugGxo7Qz2Nc0v15778/11ginM5Ro0+mFiR3e/ge8IX6ZO88N3SYHUPoXTyma++1Y4sE
imqE2WAB5PDfPExR+fnfRMQZ51edKwiYEsrznx3Fo1YW6vH0jy/LozEW
`pragma protect key_keyowner="Synplicity", key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
piLbIWVV/0eese0ZYnVGTZ5vTc6FzU2L8xPAhHPBnKw868x0sqXyhPcAH5kYILrV9kerDxnU
WLYkY/Hjmq+t5+aS2sU5flsIjtXVx+SEsAkppF9AG9sjdqm9YKKGrBiuF20TH4NttanPk6/r
GMqjnntT22wDwKvR/BwCWzv9kDer+KJnNnjgt6PuBRERAtL3UaDfIagPYeIaiyQIgccKN4au
mSStHF4uC+wn3Ux2EYYDVCRGCk6SZHYgBCVbrWEsxQWAQef9Bo1IYLeI957X1e24IaSCdpq6
kF+e4Kn9Ovrx6/2hfisbmxTEH0zj9W6Rez+2HcyIi3KMQeq9NuHgsg==
`pragma protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
Cg4U6hooni8yA8JKtB0LCsg0VmCHFH5XEGP0BmSbZy9MT2dTIHg4Oul5bHsE7LLQNgRjsRa4
0uuz8n0YYhcOh6bYk5Pa10GU/zdK6g0gyqOD7OVTD89Te/y1sTVnbHnMFX4YGWgCml2QH6Kb
/7cZQUjwCDAl9DNm4mZxa2PxGwhYSzoAGnnPPi5P6Ex1TbJGCaMUW+uRZThKLHTztGZQ9Kfq
DPfnvGF6D7coKSFBqlDvS9n91DxyIlAKdz41VnNUj8DnP8n9ZL0nAbaUR8usD4p8F2nNfmNx
S+alkTstjiqWMj7QwEU20/VahWu1IF0/VcUqDBXEmandwZIOAgr7tQ==
`pragma protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_11"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
JIQeCIHtYKUbjrE+Qck6VKUkdPuL1MrRcY/gRb4PaKZ/QadBImETH2SIDCyUDhmkd6ROzrMf
5F6d2hOPYksBupO+hEFeueHoEC/NMOLr+Q4kLdeFyselJWt6ipE60/T3FqjZeTXjMyJd47UZ
snhxwLAqxUqftKKOXhcRrBH15zLCYUbT4Hcf2fokqx4t0z4LiqYwx7zx4Pm66F91nIjN9oSY
ciLYTh/HPDHYvQKwDL6LmAqZ4FSQJZoXIHEsciqBRg7F6VPARib16lx7oIR9jAxJuJ7qq/0q
SBWdWdkVS2E9y5P9piRtQq/4ji9noH/gv+r+wiDYjOMOdRECvp9WaA==
`pragma protect key_keyowner="Xilinx", key_keyname="xilinxt_2020_08"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
OiV/DsdwhxmP4nsQKclxfMckOVs7eFfuVn2Q3HqwbfXlczA5FPuL37v/m15RUvhumUW4ha7N
EQnA5QPu+BKUd9DdSwvLYZe+/zN0NaFswaILb8FEfKZd2le8qYV2FswJTJVkAkU+xyrIeR6o
rQDcN31wQEK7jEkN5r/6ndBkxuhRw0W7KQv5Y44lymLI9uSNhMyRX3ac6kHjG/k+qTVcXRaX
OjwFsu1ZeIeX5oNF7nrilxEHmJpE1Y/RcXXE5sS9pFXoj3D6ZoDpOQYYsv9s7+o9laTPo9eA
9CnjKyOMFnatjZTHwGxieWXnQL2D3PJpNflRylRlcMEBRLfkTddLoQ==
`pragma protect key_keyowner="Xilinx", key_keyname="xilinxt_2021_01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
KaaA0rxMBmXX+3dOMTUMseqZwC9cWcHKaSnD4rYs3ui+u1ePxJFlcKv9jlB3snS5qkTEty7f
QJvo9btu6ZHYIVU2ez4w8diUKyNcY3d74PYx3QDazSRr7pUI/huDFyV/Q460LuhqY3MwEbUY
EI9+11ag0QBsJ8cAu6nLYB9VshCqnsJQWu7rKyy81pqwP01/WZqtSR8VGQl/l3XD1xgcOYgL
NcvDDhBvx9PkCgX6AJgkvtPqTV1GIh/28/2FTTdsUW6bSMezA/9xBiohhiFLgfbSTUXRWXlm
KEeOeC8fzyM1m+CVE6VD0DSaNPTDD30zWGwkmt38UzOSeZABoo34WQ==
`pragma protect key_keyowner="Xilinx", key_keyname="xilinxt_2021_07"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
K2IR3SQybasLdEcT6t6ZX5yU8N8MhfoaX1DQdXCHlqy/tCQzcByKV9aggnW59g/0mhAODtU9
GZL/ITOUEkHW00GjhdydirYRxV0mCp+06zSHQjHX1HY2PLimXzb77yJZueuuCyREjN5fhKjO
qX9RHnOu6v9ehavpA4gcOhhQ8m8w1Mm3GOKq9fAQG2CtlzlrX0/NJsNE+h37R3WVkk1bxsKP
LUPZyfjApDldh5T3nqbAuLWIC84Wos0JIHHCuRJzdD+iZEN6IDgtznkXj29ev1CEZy4HnrLO
BCWjhp2J6l8zg/KmIoDNvglj9M6ukjVoe6sUis/mLdI5Z4XgyKU6+g==
`pragma protect key_keyowner="Xilinx", key_keyname="xilinxt_2022_10"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=256)
`pragma protect key_block
v9ClB37aohYv3b4BZBA31wB/3evBk46CCwvK28ehydpV4xUR6WbzmspmwD7I7llIlz7juWam
KUqnUwcbtjuyEyr1eAQHFd+iLwzxKg/eqRxOfaMJTNC0ToW+N7sXylC4PYqSLoso4QVObLTx
ajEG7IEc2wwKDOEunq/dCir4h62yKI5gklM6Clxmp6EaavH90Xg4A+HfXok35uPfziNljtgV
T8RU5h008Jk72OhC8sKYT/L0dlbeTdZcr49Mw+gNjMDviQi7uTVzab28LPHrpVz7l8RSKAL2
xUyaXlhLb9yMFS+rlaDxj1tJOUSsvdmkKizE5usBqvd8WfojaRQM/A==
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=72, bytes=40128)
`pragma protect data_block
h5VcAA+5wfJjHMYZKXxt/yAPG5rdQwLrsfkasrAbkhgP+Am8HuYxLquAUtaPg4D6ewqNY7N7
APV0arXYgqYgmmsIDgCbqVCDIjZfjM/bxQSnPqz/su+24y2n+QmmvgszSj7ebH1378wxlENE
MKDQ66m0+pyU/reaDwQaFnEAwjFwMsSm0QPiqpbHMT/OBG5fJfl38R8quvotH+E/xlnpF6MC
5WfAgFKzdz4f6AuPgDNGbf694uFRw+NBu56TKYnPAZuCLpH1DcyFUuKnFMvGpPMKPV2q1RXw
k1hxBzpVtLKIysGCL+S6fMchLehSugP3MjMtDaav/cZUK3BCCC0nKtv1/cFF6PGYU7HJ1LkD
Ymy688qoE5b/LgX6IP75Bi3o5qLoUiKXjvALDtvE0YTgr2fGFJuZZOLGtGQgrQBxpHMrb7az
EMk+SqNeIPkjTeYa+tPlpQE03euvXHN+hlDIHmg4Aq7iz3ajDc3Wf8Xi1jK76Z/wD5Z2VAjR
dM/dHGDPHzJQI9QDf/NDXLe2JsyUJbmWC9BYt9zVI0Fngv8voXz5x+Nnft3ucqvSEPpgWuEg
mCxzxBuZUH0Wclbs8ddMCwemw3iK36hegfVYwUogtHJuFpCsB03+OZUNgy64isk6Jdg5oL2o
j3JvMPzH599gPvKvZrZyjid4gtZGEN9WzRj0YDrmYpt9khlzv7jPGTrBVCLQvJbZR3Gs7dFO
yAEa5NMb/h2XkVjjWGmqmTAXFpWsIypwg2bR7+6cVl69B4yZxCmVew3w6iuA30m7NaV7evoE
jmijaRDyl3zOoU0vc0zI5ysr/AQfp4/bZFCcp/+gSzLa9OZ7C4Xn8CH69Ev6lw/0/78mSZCd
0ugH8B3UK84XxkGLp2Ri2jU4VyPXlOMoYn8B422yAn4oMJo7ldBhNYjFxsyNxafRdqtZjCwQ
zWKuH8qxJ5e4gfZ4A1HioarsSCxDL8wg89lbUglc2cxYq7R6BaRgaIVsP7DOp8gmKz8Y5X6z
zucFB8yegrwnTaNoU4qwIG3G/tSUjsXdFbxdpTqrEKd59ylC2Ver2gOYl5tN31eF0n5tCCaC
e+KpNfMfpOtJG4N3QhVolMfaCQFt9vt8n55VJPBnhAbq86KpUNHc0bcJl5v3/M5rZVFYex9J
qu5quhu0sq4dqZiAcyDD7Sw5b33NJwFh6wBwnzq44WQTm1ZyZIgbILnUt9Sszz2NOQ/Dw/NI
hpcg7KpZZ41fh1HvvtI5NAmT8OLg0DZMHl6jc/nlSc7u+GYJxN1URoP4QN0FvwNyjKL3nUbE
USq0UZ30eJ9aSHvNJ/566MhVcpFHBpPab2ZGqpwHhdHDrEvMGCgbYrNJlIT2PbD5Y1x9kR9x
TFlGcH842RHmfjrvC5hVSXY5yxaRwYM3vshDNo0PM1vYuDX7ysIbRZXJ7DIfP4b7ka+UGi73
1p4kdYqVCsjZlljVZ3Me0YXndD8Q6ihuif8CDwNniK96hE0cJB4H/m3iydx1EyqM7yJyDVHU
TfN5Cn1HhPFF1jNkFNbgJEm5sJzK9P7qv1t+2F1u17tMQ+aY2x9aUJrVBH4ytQ/ofmjMguPw
4ru6CoSGfRyP/nJ/NWohcYuC9GzZapQfOdatMx+oHjrEV5ol5INomQuKHGz6EN/ybZJ6IK1j
gLvQNFTOC+rSsH9bQyo3AbhVZjV0lxZV7cw5ZETptHZzGnzvwM5XxDdnQlwhono+ZUNGGiBW
wfn+mqCjVH6mOJaJqiwwfyZRKMQedol72JrGJNDfrO38PF3s70MMK4tIUZiVIdn+PeU8hffh
5S+vdN4jcqu3YrdeISt/tOrDw921pTkdGG3myjIbC0o65MxYqIg8RcBSXhUJEBKvckTynQHC
FMTZ8Sejs14X7224WOsm0A8EJV3Kp2TaQ1cqqL8C0L2HQYQtca7cd8E6TLCWSSNJDAvtgED+
3k814YLwfbde+vjMMfCLmCOetjVv9nM/8VwmQQaa9BOt2r0KBhII1XuE9RQl5iBdALOtYPsB
+tOP2UePD1qJjhY/9V/3Cba5BSGTcogUV8ra2ZGoslUVGQXkjURnAKIR0+FSTRWOAKzFxmcP
yZr6Mth6p7DGGQcrEwnYpR3941qA4MPw4MK7L7Twmc2++iO7g5bYmG6MWupLUdeOa3TEmhOl
taOm/yZroy3dCqnryGBHaPtRiJirhylP3c7C8AarnLB3Amghzo8A27x+/cGhuB6uV49xpHE+
vfRKpM0eWGiW3D/J92de8Hv2DqiH9Z++sYhmMztN1qJzl/PdLTAuuiY7g+kwVRAC1hqu3Qt8
4uU/vDYn8RwpmCKKI97ZWqggmjapBQJG0cdRi8XMJPDcL6f/Jx7yYuvGq/cDDACEpgv94oFi
/9Of51J9tEFT2YUkEKbCKA+W9c+gYi0ZUV5Xzc33QOBJFbKHWYitUsdHc6QcC0lEH7GsQt5v
65UOg2jXcwuVsfzBFy/XDcskEgSyKzsze2VaAMwvYhV6qakk0qVBSXQgrWy3TGP5ESRkcn7b
CSWX8bxBwB1QCbWQiJimR25csTZNAOytv4gqRFhehCfYyRuQq6nR0V0TA06vtYKb6qxVBeLe
M1OoccHWI/gmrmHm4uodd3fAIVY9z9flD5CkgN2HG01CBlWzwj994iSgt0VIBb3pmC93sh1m
yhM35Qcyw0Yv+Dt0LafutGCzNR8BfIoRPkzmb3JBbftVDfRH53z9R0W/aWE7FmcWf0VvsOdl
eUJeRmcqkMNjIOR8vtro4xRgwFbGvxjXN6jHUuMMNcjWnaby8jV3Nr7/FTw9kdUdAhNNWlAV
mPopxaGhLsu42h8DrluhJt69wcIlLtPoorn219pAcRL+nJ7eGroBgX7gLsjywN3283qpOVGs
I7Fos/dLF3eU/mht3buh+vTnb6UXV/FTXGiaPy46gym4ccUR0/Dari2l7t52I58e3sY0ToTN
CHvN0OCUTYTTWE2pasE7e0DzWzPJos7OXPzrPU3PR08DapDUvJvifWXRS662QXrVcrokueRw
Dswnb887nRQJaj6ifEXtnjbbahqfmmYYPILHc2z48c42bU3Y3AgjWO6u9fAxO0vDV5p3KaHo
YSjS2vfiTxhjSgSJrylFc5XP7+SVGyjkMLzjfGDv4lWawpwIeavMEG4VwocR/Y6GzkvIl9I5
+eTf2/vMh5jfs6jEIYhmFEL99HSPTCki9o7rBdOndoV108q0toPw27PNGrf5cXOY4uEGpZJz
jjtp7Vf+qMkzi/quRYXOM4CVvB9cXUE+A6jrhfEqlJg0tw6WWPKuGZHUTkQ55N78Zr5EZ1vm
mvJeqcd6jlDOFPAILMR3wPSKxrG9cjW9QXlQOdcoTvGgpLRG/YfQixrIud6FXqsa5sVgDd+R
P52QFs6KM4pPjHKgHuM53LYfnVTyUpmNvkX7e07QD0WdwlHfAI6CujD0IXxwo23OUrOBfa1z
QuTV2aRUmGlLyeb37osAlm1cTYg/Um6Vh2qzMNJJpXsk2mSnu/egHSPB0TKM/Xq4Smtkj2RF
ug20ACGRJGQYwseS8ygLyNYQOVZtjALjgcdFNpNX9U+nE5VURJr9ESYvpcUu8FSPdjjSexiQ
jcxqtVV4A37JU0YKrbwnWFfCjFw8OXy7zPZ1MsQMEP4G2JCazB+Zfbd7y2+0nWErHDJoLS2O
PosiGy0DjNkuFR7tFBK1lHvQsPrGFfp53O5wkFaen3mP0E8kHCMLK9qvHS1UhEXBVexT44hB
HoggO0BxNXa5HjVRUXfgbEhgmdo1dTgsYjLXZT6Fkm16rElo2u+pXAo0L2QJ/Tktk9YspUEQ
JOPHNK0hQG0DePsI1DpH/l1pJTaFoZwFw1mREwAW9iTnjprGpjgaLoCune1ZJEA2DtDo9pco
TOhGWafV0le8cfJJdepwWb+kKNwNBP9S9QKHJtr/lr0GuXB7wo0v8/bw314xTdhfaUPfLRBu
OYhuqQYOvWt1pPX6++0Vzxsrld56I3C9Mx3bDyPOmpmLV4l8CNouhIx6U39DPiwCJpQLXfGi
/pQH+GqrQN00tEP8Zma6+PzAKpOODuL0NKf5E3kD63LimacKxtB4GjCuW62aiVgzIiI5CPdP
bfzJu3pCdLfT3LOUQte88+Ij/caX6FznWjeHYdM9lP9peA8s2ea8+PJ9SiG+GuAVRfd1fqzF
OD1liV9OEnLTwMRBdtWp1aYUKQ6PgEJ5JkZFMKf81zs3w2sxb2W4zEMjSa2DHF1vSBX6EFUA
y2fZbvKT21NZfERiAWocTMUcrOGzXni0PMoR/bNRa261Uki+oQkviIlxpACdpVWUOzVh3T1u
I4vS2wKlmp9uQXscutnwOsOZB/nM5hHm6wmObVuj/mBzReq1dlHnFAZvi5wIPXwzs7+4/XQ7
X0KdP0a6iI4lmbCMcR2A3OiSFfbgjflUyK15b33Vegqk52V1fyWPvHnT/WU2Wzg9J/HDcbXY
Mp7KGB21PwBlDCHBncUGbt2hnhD2GHRHrjyyNobw+/TqEHzJSDnckWIRDSQ41o5S39YE7+h/
dFO8kr734lCdEsiFxLtpSa0K5ltGGTp+ZJZMN98f54dr/idiEPVX3vnj4u5sHW0BzdSTqGeT
L1T+H42csRnQnd3R+2ErK0FWzNLLF5oPQAzT/UEa5SBYQzWZugrvrUblzlrNu1XO3LwEvvdg
2GeIzNElAMC63Sc3TVXmetPcWyTR40H4CstnY0ZNsZiwGCjh5/BP9u9iupzZ4iy3DeC/Gpb8
jNlOvu/xqlVJeEEdlx2giqGMQaEhcqu0F7Cl5//TjCjKk9D7uPWsQnqmPUiw/u70v7lTwB6n
UAr1Yf8Eg3FrcdMJmN7XQ2lPvgSOHzgEs31MGh74k0zrMgKLbrryNsqfHSau5UOVsau7CVMe
6ZaphioK9c6NRJ0HqipKnCOBiOhuN3egtwKbUkt2Wnm9qkh9OYtkkG30L0aak9c88Wp0dMyH
cxNI8+2n3IT/3GXCnBV9i7K13cuETHDxtyaTti5DIpaicu+B62jyFe5TdS+ZJ27dL07Bq38r
4b6VBR6POXL1BWDA/jFYfxwGPLucWGh8NYefifKqEp/hTOoPazaYGJiQD77UJ+UwixAinN1D
1uBRPatvP6AEsvmmnl4qv29uXYAejSoJW4hN4eqyVsy+3qdlW4yTL3J80XxB1jDKf1+ZdSdS
6ugjRXjHpy1KEcy+00ObWlgykHv4XZeGCUkUN3njVmUObut2uSSX+9d3NJRc1infywUR9Vx1
gbEhic8L/TZJjU3OiALcOxHLxPSVuFS0uxKqH1SghSadY/HeZSnBhKCDAi7odvMFQT+p2njJ
H9n+5OeEYs8dkPcwiUz1QrU8x0exaB4jNr58bdvNQd1HMJYIItKWqNObkN1QL8ncs//KQ7v5
CUHuGMtyZvEIt+YeMuNLmGlwv09zeOHNZRC62BmKmOglbO+O9350H3nYE1nuk1tuGVoal/dF
tcu/pwXwjHnAETmVLme6CjS/lyTXGsiIkNmdH2UTSkhqrxh7teNsc9TA0yH5M8yQMgpFRs0A
E288v9BNpRpL5lWA611vQ7NbH9DvZNuUNnfXKk1ENUGNJzdyrT4KaSvERYuLQB+D2PjWTWcq
z1HhqablRLXiDjBCdp6qhBGXjS/twPlzF/uzoBqV2l04hlCgG6rl7Wk4qWxZN5+re4wyI7RP
8znj1VLbgmqzEJ4mxmjhixPaY5Gy59ujKny9ApaNRj1yOHfH6hdSuKlx26ifOqquEQiKzDjk
tI2KGPgeufITfrJxzMN8YdQkTl2uBnpOTrUN7Ubu06hNrZu8hfh2lV0SMaIJQQXTlWwrbHKc
4AqHZf3iGO8R1gx6ohkeoelse1vuL3WAooTphbqiXR3jj5zoqOGilbkz9GLvelOxiaHq2iwN
GHc3BJIgLEsRyMOjzxrMzFWEcaBdrU2bRzgzHWL/1xnrThGhonmzqd46FzUXkEGFLZPQApEO
fTGysws/yzkS3bKLJPG+sr2OWHQrLpSei0XJ3Fm4AH1WR4ys7rl8rpEcChapmZkNkI4uRLDn
LZkWtamXpP+P/dRrx+kAEr4Ya4pxaRjYx/MQQVp1eK+A95dmtzxOkIQqkC0Uf53/yGk8Mw/R
rbdtRRnZbeV98QbcVQavCBxIo4lwSp1EvIYhqOrf/09XCP3tUpOT7bKNuMpv3sLbFKCNOl6J
EFMPU2goP0aRBErsAzrXkq47xQX5p1oPtiLRRs/d0VEYN1UjifZv7lknxA6ZCMKcy99MQLGG
yy6/uxNXjaMC0fRDaUrBljVmGEZ9OmWGnE+NMiSpMcaH4Lbq6gy6pn5nDNJ1hwH1EhBgDlYM
JnKFsS4J6l8xDYSNOB6pb1hyfcy8IdoZ/mtNhbCMb9Z+pHOKZtlrHpIJC4qD/VaJcfQkqPWS
KtOHoSmdvBUxbjycf+zfwPsaniwDdGoAANBtswV2FqrXfn3W6oy63PcIQccWx5xQEJhTAEyH
Lb2CXoWQO7stLtI6888ovQGRngf20e6TsHuyL8yuFwdXbO7qlcoEyMxivpRfyZH81/zDrWNk
AFtmX+f7bj1HiiueUepGgc5+XUVUDytMuhuPnzTr182lDNobhSxt1yO6YE0qi+On3KlCX9Jt
81DShC5BaGvf+7DOBHPT/EUH9z8Gp0JXGR5faZQv7sePovDUL7c116XdatB6pUHUSPF7WDEg
uugiMyM8rH5TvqSxKqktZx6YbXCe+4Kesg+EbjzvpIpK+E9weXIx9X9/A4aVeyosE6JKl8KA
6uVWQCLYs4676L4opvZAG8JFSa52BUZG/eW4KMq+ooqGsKC/PDagGaa/lutatGNMJBssnueK
hrMQZ6ama/fNTgxVcvSZOvxV7qHwfvG/iCJEbH4L1gizVIp5rV2KfUqhFGsdZvZ9SzdaQONz
Y3rwvDHzauOFjcz+PtEA4xLsUT2hHTyg8T/O4XLTelTiy9WgHMLwtteZdw69W31KVjdvpGxs
bnt3Ir0aMy5t3khe8FPoC2AI4iik7cnq46rLVYKAKC31VDtNSLMNux8taMQnP/nnIRW0C5Mi
BSlHFT4kK2hKYmRfQnh2wYFDuqEbmGoot8gfMs9GGarOS0JOUinoNwAg1A0Wlyr8Srv3iQ5b
B2goG+ZdLy7h/Tr5P5DI4QscPcU/YsR/AydVJI8Xjdze4lgupBddv/o0GOh35Qgl/E27+9Db
CBsS9sor3PSqtOZquKiJDCcG6VGNalOhQQGSZdwuAGrrf7r9zcQzIWLPOMY5tZIA1NuZii3a
YEG4XcR8tHLuW+J/rrhvz5NTC9yr/K9daV6f/FCJJ44f8LL02bLXzm0PTwf/CHkRu1AMEkMU
DBdGCYskz5S2S0qRLngqu1pj9cQ1cumShL32mXp1DkFv2cuGT8vXvHxsBIrFNnxVcZ9oVeHW
SriQRfDqFWTpGfXOhVHXssjMf/n7CBC6X0ngPlA+LFLT4oojKThNQMdxfyYxPFKqMMSXr/ot
MeUe2zyGpEqiylDoyQq+YIz+3XbRQBAAq9/kL4TzReAJQSJnj5i5C6YEEc155Y/wYe8sAM2X
ZbK6+xinaQxhrgBBvTkOCPMCiLRmViqDXc46zdpGJBzqdhc3RnHP3cev/C1AYhTpcJaTGTbw
348puDX20fc8zQxzQMAae5PVd98gk1qNFqxVHBz575dJKb3B6qq7xRltrDKQuC2BzTZFd7W0
LoVIocA2n7I8ywsKT8QRwEzkybwGwQI46sU5VLyS81vMoi2aStbSQoPngzuZXiwNv9hnNfax
mnWdzhWqIJzuyAi0zcYONdSIqTX1Eu0dAb889trwM9cOjaRtWvyjBW6RUoc9e4AmH2zCsxdR
3++L2rC4j/vQHljNKoZm7wN0Ke2NvLz2j3YEJobveZLOOl60c+NHbdUwc3HaPsgUo3qVwNvs
CN5ix4duVRCRGgBy60WQjlO/Esh3MJ4y5oe3MvG+DA4H2hHKusmZX3J0TzgYpYnMJgoUIOzt
B6AL/VghbKhpIeMJM4L1BA7PQqQqbSz9dqJiyABXqUeG3QMegWGJ7TUCAHiSEU8qDhkqPNfl
qaQNY5b1IDCesdCLYeBlZamLCp7Uar76zIcSP9/UDSzTfVr/YbkeI0oEc8kXksGORCM58lbe
cxsskWCjdOY5MM/os48CR7KlqtJfMMPsuegy73irjgbpueaS+syuGsS6An4YoIXyd29RyS2A
c/j3P+TVBO22cjjAC9hI2dT+kP2wcwFuhUPoyf5wtAxbpPt50nmPWTzt5MHtmjtQCmCDnPnh
D1uOqfrzGPYVGwX/8qfnwo95m/YQP42LVf7JAekbvcI3/Iht/cfr7b0FLEctGv5Q34/RQ+VE
I683lQsRhFY3GvIm91KC0Ok4sdYUVeShcjJT718ZMMUtprIz7lhUh9F8GmQbBhgk5Oy73Vle
sxdReVBmBocHzY6jnzdgqdmhUDex5+s7TW7Lt8/i6kKJQsxOTGvbZV24F1eBGL8Ej8Qz3k/7
5kuwxfc8C++4EVDrsnwW4ymdP+2+kzEGVKQBTgLb4kRIVAMuPCJJkkSTn1WoslqgIptr5Nme
1/EWuPkHqYh6Dj4h0MXPHU7dNzzdzg8caNY9YyJdMHM0QlqEDuQRzoZo0jAVo5KxRSgrjO//
LvsHCvxpoz1wGepnbucaL98/4uBp9uwueLUjj1SMs72z/gFLdh8L47OgLbOt1oV//EUQTXqT
EwpnKegmflY1+tT0k9fwB0VxTXRNXI0le1wkYCZ1Cjq8szOiK2us0dzRpY5z83A6Se6Q1Oyl
ZdxI8Po6y5c0rtpaayxmTUnO6Uchiq4FUeCPADsrnYZy4O0m6OIgBxsFP44ks1NRJBYX3gus
8kZe4JiUR0OjgH4rjrf8Sd7t8mfJVijn8nnC4xJ7B71OZZcsqiXUgaibIzTGaN1JhbXsoa91
G3/uYq0Wq6dbvwximJYkSU2FK18jV75TsKVrKgHr98pPFmbUtInw9HhKdwg+CSkGRIEOtwOd
N0W+N0Z/Kj2JRln3FdXxyVBJNLCoHa2wxC6GTCvkr4IxI9gSyiHZ11OgrFNsRNn+WcVjiuns
PYna2u4Xw+2aSGZOfcwONFftlfF/jRDcromnPbnDS/TzPkDwNhMOjhxbkPKFvAS1xL3qi5Lx
z1sZQQSg5UQncKqZPrceYTM2GEBcXzcsWt7GWuAU0rXG/RrrGlioPV3fdXxeiLUeULMV/30W
J/vQ5yyemv4CW5q/+rzJRMTIkTGMlSV+9XWs9aS3wzZSqlz+WqiTM7AW6WoGoHx2JCHoQYDn
AGA3qI8afiuuUwRHiqp9Btb2RbQcNfN3dMjWD5G8QDwSx2KVvR7zJTC3e91lF0OkjMxr8Frr
tLpzeEDuthqJmmKS/8wTd1VK5OdUQ1SF7/UBVgdedxT/Do84yO/47Ooi+xn+8BPV/RptxWzP
GYez0xck6ylW74TaalJneBYcEnkVOkpbdM5GkNtazNfXKbrQWfiT3EESgTzP/YMv4UzUdBO3
94wP49pUuVcLHYSyfZUkRLVCIqX8EDi4xXfFKOkZLD/pduJfvw6W1jFwWhqzZrkRIrT6heL8
unBxuLeDAkKX2yCh+9kT9Muyv5JwgnAT6A9O0x4VXgd/Eq9kvxUcdKEOgaPXhgXrlX5EJz7+
VCsrY0xqhYXGzmCbi96zJpqZ9ucCek0c3aMO7uo1MuSKaDOKg11tSmlPLcNcfSxuG8EbrhPx
Icpy8LFaLrjl8T/l8n8moTGkR3UYOb+3w3nic+mwE6VP4SQXdMBPOVzKTLPUgkOF9kcWgbdk
jF3oFbVV7uVNFpEAxoSZSWfTc/4Kmn2mc0RXF6voQ/osyOAC/U4k4IjIIZK1fz4Sw/t27LmH
pS+302d51+9Ddy0Faonaly4dyyeJbS8VTlVpl3mmcBnikrnIymUBKZ+8KFR87HGuIgIGMa1o
mliNlA13EcHdymGeAe2ILbMWJP779wOg13oLQzkQtPFIo9TuaeSTnU929BsHPK0DnXOcWptF
BeU37TofmYBBXiGM2bX0HMF5dZEF2uJxZeJB26A+6iFfjSz0ZJZQD+UWK6K7mJuk4R9v1ufh
598DntOX8wBYJq/GpMPfR/Re27TtLatVHvcxfWw/YCYtUer39p9bZMg1E4AZBzosrOCsYXBy
0d8bu64AL4jO1sFNNNL+eB7La6UmmYUa7tkdg4nhwCeC1aQlV/PVEzbihfgNpPPopgcLhljc
e6thp96KBwVKX6l6rVZLCTsUQF6ttmu9ZMKQAQqO4Jh2tYUN0yC2CSpAyfAFk7ECzZRQCwcz
tNC+MmkXvCTmDDBsyUg2pXdWJ0OnxKwSc5t3Hc1gZ542UI5F/CaWKg9dhzhePMWHfO7Z/i7G
1Kditesdmd3q4hpUzbOB4J7ehtXnjtFBcn6G3zfLgayqbRuIm4bb/ogrrZaFsyIV73xK7F/d
hRkE2IMrg98GKNnPea2nMA62ykfApsuf2IXZ+CIgrkrpyVEWTg494LNAUQdehvi4JXKA0OA1
04+fHBCfaBI6r40FOpjrsfeVDbWRAgfIkqqYq34uilDxn5ahIyfdstytZwAKTiXyQrOL8MU9
tgkDOGC6DXX6RBBWCrFLt77BqKd3uwI+pCVhD+Cmasmk71P70qlvqSnoOTOrniWQsjh7NgpS
Oc4794IXW7FKealuKOS5MIu1SJx6f/54bCb4eHI3tcpf0/BjswhDWBflLBTuvLVAX7Rknxwp
oaItk90hRTUNtDdk3Z+Ai9xDME8anvGEXyn3PMfFbgZ/ROobSmsyHD8g0s8EQT7j/p4SfMNA
bIRCwXL/583ifpCjKPiQwhRttvTmiBmSpCAnPBQVQZRdvDhA2RBPSexMlC4l+ZAuERJ7iLx3
EnbFQAoaE0Rxc/oRJijY+yTEZbJqL93CBdV3Y4BqjysMOjFpDivyLQqCp/ShtDowflJyoAWF
Zn4ACvCRytP+xFZ8qQcE7Yqbm825c1C1WZTNRXmh0vzBMx1hIK6DOkkg6Yj8czwGF+CWfPQY
rmkD4utjv40wvKRilRXvpSgrIVq0DktJhk4obszzSBM/s8RXErmFo6OddRB4Okaiyf76xabL
OhRqKEJsN6Msx4NacXNlJ7Mo5SNTrSPf2ie4M2BUuh/xXrkK1f/rfLH7hBNAea7fy1D+XrDF
gY51JUvtqIYWT4ux4kDDMf3nSm1kRYMIUWscicA8Gotpq/k4WJtqubi/MFOIAyBtYGSwdGKs
Skgw8fclBU3wc4nsSf0XCGY/HvH+GDDTHkfhURtiCkSJNxH/CpLTY4t/aDCF8CXpo5ag7IBx
P2jB6yoTP8nVk1QEk38KAGrFMxRTIOB07fLOT3Tp2661In/Off8gXBpBQ5/t4AyQ3YZ/woNp
xjU49FeFs6F6gZnpkqvVRWVhO6QodCMo2ZLSD78QTNLwBvAQCWfrHk5jsdNOz3E0EPHIPMSj
ATk8MJrfPoGouwkUWufKrev23qt7GEPNnsUAenCgzraH6hoCDzTO3vYg8HNP7llbHuQCHYUn
2SvKC+TmJLrvxCg12qT1N8NGtNT45pc7fTgJtMjMM4lquxZqMJB4nIFJGJDHFn8RL7ozBEd5
vTCASBwNKVSgCmCGNoQpEqOUis+r19evOnhkiJ7bp4KN2LiBNC9wTUKcMiH5+Pb1+8UTBq2b
JKiS2OWLLXr96U7esWoS5vlG3RKVo45GwXnT69wcLtulopAKssPN6cOGuIHqEzu2YRo3QidQ
9qraZvHvfxSIpaU1qFnM2v/0zq/Tyv3PHCRTKdEo79ecnV3xfF40C3JaZbXszw7Wiz7aczpz
OmoL0W6848jMWpzUswE4xoAU4EEPLf91ejYYoevoYuheGGCP0hw08j/vx26z6ALWPXHdpOPG
O/gKhS940/Hz4t0q24QsShQAaQ7x94vJo118vt9XVS+yTtRs/ndaM1WwuHIa45bOrc8UlnZQ
99aWiZ8TgfREzk9my6lDt0XN+MCxUq5de97q42sPnsM65HnkTJvE4sDBB2R4Vexju9o1bvj1
/e26rwjVxXev1nZdYhkDbYoume2oSEH303o3LRIG4GICmrXYdRBe9fvVRbbQnZ+4PoP3jTTo
aN19agyvPkneM+jv7wql3347uFVE3hFn5vGi3EHmbp6v+Cgajfom8inVU7s5CqlidIVp+XKV
byjx/tLHIObqpkY2VW5scgvZUO7XXUFZoCLpnGnbRPtAdFTLtfAdyHH4lax2+wCeuXtqQXwv
WX4ebQsYC4zOWmW7dVY2X8Wp3kMr4kwDbOx73f4HMZM7ypIzO44w6aqw4ssHXiWv8KVd4Xfv
CGh6qkTW08MbYYLoX3zWH3Mc8ISEjI2l+uMujbaWuRtgNfKQAzs6PCtsbwaG5SyrNfXUv4Ug
p88UtD0GbEeWDVRzCGUM8H81gJBg9ZeZF7QDmwvdTJKegRaaVzU2HRbrLq/d59ovwlNAfDBN
uyOgSvg0XfLEnsI9EBB5s+H+gMCaSguEUkFpTgfX8R4+m/bza/alWun22Q+38CnUCDGrg0yE
6xFjsb7jLTq2uExTnNfPnRtoTkh1yfXuF2AeUnYDdsxtZ5BSyCpGAhlBotABKEYzfZdEr4SQ
K9i1YP7uCGqSdF0k1iSxnf0CabjAWnWjo63eySUh+sX5aqUy3VvIU91vLyj8zWX8yt6IHb2a
gBBXQmcqQEaFOGmvJbqvFv36iktdLrHgWbQZpeSVjh/LtFquzIDr03faWQxS6Uy6X5BuGKGE
ZtfsNK3VJ/UNPPGE4UDIpUL9Ym2gpL2wVuHsNIjHwv4b40vAoMi8pj3mfZyiIWMq2lGMQJmS
ziKddAxcpJATk1sgcbv9Lvs8UCdzcvnmCP1LHn8uxoYB6dawayj9onjyk6x7zVHNVCzdFEJe
/Umsj8QZEUquIZ6tf3zJI31QPB0iA+0jr6U2CaVg3BU2t4O4yT0nM2UyU8sDFQRngbgyz8/R
lRI/P+/T1ticXZG3nEg3/z8pPDPsizbdAl5KITJl25fkX7zS9fGQSJSBuxMGFwQtKDuHAPw9
inrkWgQ/tVdW6xJM7jm/Qlm8NUUMUIrefsZAN5MN0TKzYM9L1Vg7YPNOMjYjpg38mXyoxerV
KrAG/bLIuC12dQF8BxyLauvFsva7uz+da8ThElPt91PIqjhk/gG/rLxEixgwE87qjSIoM8o7
y5lInKdpUTb6TqBoICDP7Vns8QYaKQDD+xEZmFm5mlhYW3NDBSND/XHElz/ShYl6s+HwRm/o
GBCcsGFt3sy9He+1ChhKTsSvx9bsDPT3jYIl1iT7rZWvBUvlvsrgVg5xpUIalAKurTXJII1q
uu0pFCwDEmxOQLnvusJsR1RUp//2sYmCpfxZhHcG+0ZcADEBnh+kXRvYN3Y521wz++UAO7rM
bDlAJKVw27RatQtzMvo9Z115lGPaxXlDl3TCXY5qK8SmehpoLi6gsDxIo/BvBEaYaXKiYLP+
xIbXPY7gl2ytgHGQKdiK2++at7CXRxW9AvpnuLqTJ7D77Fijm2NU0dVJsNbGzuhEAw236q6Y
y+6NhKCKCOF1tvgFWQktYxBvsZqR7UZdCgr8k1wdE8cxwcCFGx/Ewj2C4IlWI0YD2cf6Hjn7
RZ22o1emteRWx+Y/l8oyLpL97a/kzfZrVYLGpub7DyU4JnreEvDxH5io0ZDXIJ+++OZC2uP1
RbgGk4iGXU8hbU6/7EWwT1u2k6MbDK5zcXtAurrQEPOLytKIQifC3aYtcX+lDE7zRvY9tnW7
Z47Z/1EHpnvwD1Kt54GfaZ83FD35Ow/+u0MEkFkP4s/qy9Rn5DuZs/Axq3glkOqnlPVifjhl
XOMykBuQfYl6tuLI0sdgy72G2PivRVT4rifo0oecHNYEVLDzVgulU21SIEFKHUF4cXq+CQ0M
HDpKKRVEH+643v6IBDC5giAzq6K5QamvRYmXSXyLIjAYJSQ0EBlALxbR233g2h+ysRtSN3qE
1fwNIIjn9ma2mOxlqkRQlOjspqrObMjvIwyPnOWGHkpOOacpoxNMROxUK5yklCMxjPAqJBko
/2LCklzC8colcDWu0thBBNUnILFzt1XyQMudEJUvbbQ9Yv4EiZkqnXZ18PQLamXVBHx3TaZd
Q4Ocb+4YNl8TK20kvQIcm/8Px8879RIRAqB+TltTd09idzTUeO0aAzim2LNvmhN0/95IZsP+
0fKW7BpidePzGcc9rsmMXrKemJxB1tSxkqZCfwpaaPs2iPkiWR07wMPq0wdlnVoLNH3d/oc/
z6/zWo2czp2S9rIRz1Mim3MqlcgXv+skDOlpFIEIaPYIYxr1t4S453xyvL+LISAt3CF+XE3W
F7l0UAbCWtw5irmvY7jyDQrKNMA9ogzjxvDzZAY6yKlJNQfOpzsOWG9UlKn2OdnUXtnf9LzY
74i9B8yptUiOWeH6A5Aj+H/AAM+te9kitJOXq9+BsuR0//tUAmp50Hc/te7S4Ug9pvnDdViS
yFKlOEK2rz+soI8QB62cuXSx+teWLExvbSkTJ6HE6x0ibSSJ9MuYwNO2KyzabhxhEVl96HF0
W4ubRcHPKC07WJkSyUh8UEC3RlGXJ7j8Y7A+WGXGmLQgYyn5Xz8vD9/y+Yyl8HkhyezM/ACj
/PuPvBjgZmv3qc4SnwzMHEWjFYRvwH/U5yA6J8LbDGwrVtXwFP8Hr6u4q5HIDpo9kMHJ437o
XnbJczMkVpx9rb5vxuYTagRRZNBRbm2mYE2Yn5X++bnivX9Q19LHG3F3xtn3CvAwdsp3yR3Q
J6f3h6mjWNaSi6S7qRo23ZoeYuwG4QAm+xGX9kt8nXJ1CorLtVCQdTw9/E9IXPnxshYZ72rL
yCZZ8vbtw4k7+IxCAe8kslIP3OmmYOJKAf4zZaFSjMkb5H5qZBniv8wq4ApOZ6tAtCOYB6ce
jx4u8f9EoAAu0y57NxKHuNxYvLC0LPuqH/pejoWDVFycEbM2nlQTvCGT4JyyVqXsxmRj6scB
OgP9XMCHGfc57AuiWKsIjAZl37UONiID3HZAjBT1m4AjhmAc/fgc/lJ/MUHAwHtFFbE3kCfM
susOKs0RswVnjKnfU7PcPTomcLIgUGPVpOAj1XX7m0N3dqiwN9pteBrfWh7a7AwmVBJRlgcR
lLm3kf/jhGsmey8og445k5Lqc/G3pBV3e9NqvSXvQzKt+xDtOJk0bvMApP5OLltxd6rd0WI/
ZYyoX8DS7ZL8qR3Q7lEsalWEA+/i186KvT4Kr59qlIxe6hM8e8WBrtJX+Bmd6GqdOEseWMhU
NLJb08qbo14igb4FFpwu8L+rM+T/7SvcssCiDTu2rBCOJW7lOFaynAzHKWEBbcTVmUF0RL9W
OZloo21ECw9rHnE2dnEkEtSp7OcWO9EpfZNCSX8Qx+rEr6SVVA+c1eMXXG61IWZpqBip++b3
JVyyRcVpTaNct4NpYV+5YugVMcRj4m+A6wfctW2mtPdIA5VfhOq2RRGk4IcihiuoDLOIMM56
x1NDOi99TnjZnTieziWTmBET/uETmVylfPdo9cDlTJBNz2cHSnk/D9Wg8Vb+W/rSd/d++k22
r5kCqIlIJdkQ7y8d16GIyW/8zY4/FHJv++D/g5i4B0sdp70wbolBx+fuVmptX0swTmpgWKKP
cdrw8vBAH0LYss0p3MCpZn6Wrz0sHfMnm1s0bI0eJ/UxyXVIbC0z8Fj9B9NxKcrrv7bVf+rd
eKvb/1zxWTZI4CxfASoJp0qAXd6hlgN1TX8byQiOhJ+EQHETJKsY1FquDh7vgs1pjgVKhINA
wOWjSEzkiDuCgwcdhqKy8VAvuPMJHd8nL1SXAPUJlheQ1GTwTq4ycfOOV4BNrcm4GFskDm48
iDjYRzYEV1TTACPZDQe6g3JN8oG/OH71DuyfXZWNyxy0wR0qOQihPTZ9hugyS0N7BEc6ilEK
4pLUxA+KW3GQV10M0YiQkXpGlNLgK7MgISDwfJINFHoAwIdZv85xJYHM/cu4lUJ2FC5QqDdN
ewHEtr39o/D2XEwp9xUvJ7NmllQSpwgIppd/oSYA0KolCUqWZqsewhjnlUhNpvikpEoEU6FK
gRxES2P4C97KOnl+wQHNmzXUi0zKKhcyqsiEIx06hwiRCVxCBiUOSQ0EFe9tRMVe+L/H1+o3
L4kYhh26isGtdDJOpJfXbTaY6Yi5BSE/zc/OEdxu+4Jvq2IPsXxgRgg0QdSdP5VWN862HXQq
9OhNT7sct/Mo2kmHO5vC7yZzzdgmVPTu7zA3K0z58/216bg5C/vt15pabvJ36RsCDZqRU1/Q
mm2EMCyfQu3lhrRI/mj+E74Ei5QYJTIjG1TMlZV5kToH3idA33uwfe0/zJTuR8lZA0Ub9+it
zPmPn3JNYJkPmznf6c99PqWvRMR+TOHECyn8W2X3NCNLzejwFRltl8StyM/45butY/QgEBW/
7PA3jT8UebgoNSZoHaZn249WDzuP/QgWTTOlhckrY+VGYnuFoL7kDt57KFTViW3NKf2/BrTD
oitTw+JC8ySCakPKugP0raG83ZFEy/xik/9UGKk+B6yvAUpejh6RnSGhkogZx2b5NfD0vjwg
dHCuG64C4YOazQXUGUM1Kr7qu0MUXtFGwoQF90vzXRnYHH34fE3cIacDUj730iDTSdXYRUvt
jaA70yoVtn3osTaCE0qepxW0iFsNvtmpP36wyYrryMMlZv3wTGFidXC8vhOQ6JH94ajtQGT3
zrxVeMRw4+LWA11KhkliKHSan4HRlROrFEF7lDU0Il2vL3SohRHWkKKJwfZuEsbPSZd9cb9K
8MdXhHS3hnT+ATwCr/7JxDFgsV2jCFiymWG6QzFofPxQOmLu/OQ6FXDTExqC+7vl7ob5o++d
hf1Chp7SI4SYo50TI8W74Xs9rHvZbXG+IoBrWEHYU5qWMNVnWoo7XuPFmaPEx/00vZrY5UHh
OcMsotnKLBLUl0opy8FtHm4HgPXAYSqsV8UA/1vWN22pGdPTh4e0RsxLqHera1Gp0w/kWa1P
nn4Hba1ApM0E70nrzrkWyx9voIWHaBYuSaM+szTFw4uu6yN0In/DicwSchUTZxO8+E/TIzgS
IomnU0mHuCy2LWGZ5avT7zSWPGxh49Ip9pJaBP9f8Wi9QMJhjVvq2rU4SGlz5ocNQ87LY2we
KrKk+eN0F/zp2xcCqnPugjsLwFn/TMaOIDQjYIlJkcVjV+v4gTKlxOxBC9WDVPNEIsw0wyNP
Novoexuo2vLfRXJx2XFWoXcdkuJq+G+76n1XOxNH4kgqXuJRohZNbk9CwMMBvobYWH72ohiR
6LuLpEjBDBh/AfLCV1E6pbROKib1fhKevamEyvdna+8Or/XohFAcIfbIuaoBDrlS+iE/1Fo4
svWmAX87lRG8C8G8ud3TteaoTEWMtjQq8A2KW/bPxpnh9OVwaSsB0HhvrVJe2n9KHnGkYTvj
mlzsUQlSJg21Osvud0Nobqkd9AsViB6HjYpK7Oeud8Xe+SloipkPVoR/etg+Gz8NK2WF6RwJ
2P+swachB/IDFDzm0Vmcg9ZmMWk9n9eyVRJ0CM6Xij28IIcVKtlfCzrfexYBen/N+D1x8iWl
Vb36a+SkrPazNmKBDWrLkyeYM3gbaMEogNKTSibzNg135sd9rxNGq+qcRiZp1cFxdAEzakaG
GF95o6TsJ3IScBLwOP253EsAAG3cLzZkPCrsGqznmz0BbFiVaNB9ujR7uBXz/8DHw3e2mrFZ
Fe/FztMws04fCIAlbEbYurM5cGEYpXVw7JFrYgV+utX3ElAnKjSUTTCstM7lYk6DsTfLU/bS
yQq8gTVS3eB5KJ/s3H94zKiQ+lg3Dkoumjjr5E6ZuKgFMEf1gSAjSdY2KQIhylxYPVHyBMSY
e624/d1CGRnsXUtkc5XDcU+HpF08OwdhhzlcJyArlJsTCiIO+DOzrwnsxkii8SFtX7Fy9HhO
r2nOJkql8iy8E5SpT6NTCnf+FyaVM+ztCmJxBHWn7bywDWHsmW/JxkRdZ0SVIZu869y/jtex
4FwumBuC3+dlmL/izuI/zl1hwH11cAjocbwZHXef/CtmRGMCztI2HBL2naD3k7MSCZUXmSmx
mWWLlAV30fAY9yRo5k8Y39gl2xcAjZbGwH9zNK6FfmzXpWj0TSwo6VUfSRA99lYPYOm6V7FL
INGkvBrELRw0kfXDnpnSk3znuHFgYq/bs53LW/aHSKuE8hn7WVcv0UDqQwMif1C7idkmG7X0
HBfQEIwtX3BHKFGZeIj36iAYieZMmVXxHyjhGW5hZzWi4+ZooaVRMo+gR1TDm3H3hwf/EMr3
qUImRRk9lWjtq3V6AeCzM6Alqf2b2F7cJFmPW7kT3itrCZKzV3H/wOEgbqdisWyQ0mtk6K0O
xOhzq+Lsf6vzBGlCYuPguJdE/5J29ECNkDNzUpMX36sBdxblVpzizS7aAtZOwRj6HbEiB3Zy
s91EhnhhHUsV8D5KHUXZOwYxs6iSnhy/qhDG4l3t1t8+g7wmKgb8bXepBqw1fSMofA290bL/
JDQAC5991KspcszvdRrj3QEQN947VthTNLY5PExCyMlTcMMOOMUSwnlph0etTGoXLcaHBycn
TxV8EjsXllriMzN66Z7JJ6wQIrY6Dmwnkpsxt4lq5p+EzYO0mQx2CpQwpJ0+9GCjDEp26yPb
pR+jep7A0fUoeXR2Ls4F6lMWcWJTmVOEjk5puqmEO6ysSLmqMob3VKtRQd6ThtFF6w+B7x30
AFFZMB+RmpgJZeeWoCdg4J5jPycH1KcNYnJ1V8a4HOodDuoUQjDA2+YKZcxrUZEsxSzEa+Mg
E2AcTUM0gtEvF1wYisOvcqj2dHYYs46fveDVIgRJKYaQ7LfubLhBVxESvfKBiU/g8NfTL0ut
PjKIwAWcR9BPCJhgWAnCASH+CJdWXiYHM194m5yNdJlbfv+teEBEpYzWV+vht80wjNBBcRry
Qf6sNl6A7si1lv6ydOQSKImzeVR+Y6q8nq4VEtweqFg9i/Zi+l8bDacARxLftqpz/KRzMdeO
ogvl5sj5UWiqSWv82M+YTqq7K9XSMVD2mfOLupC9MYoXr+9vfG2sDTJgAtaUeIMClkpGVB99
Vh9sNpARphZdm45szc8z86E1hlg84yC57w0tTZJBOKP55MSQOZBtIUn4ahFGhkaDb7DB4mjT
snincSndPuRMt3dx9yR0zxxuKUt9v/Gb8w80lE/m52OybQmnAla5z0rmmQ842qzpAj66C4UD
2I+i7njEDsZO1S3wSA+m2PIjH+qy5eS4mCKDgzkzgMPnBLRSGE9xuU50XH0m+KYuXExcQk/b
wOoz4OSKnGU3S+4rgeFZvh/tJ8hzgbo6Svuob1sUfeo2oQKiqvMA4kPKDSZ6dlgkYHolRhrE
zEx7lup+BWsIHhxDYp29szXEtMDUk+EX8hvKSqetz+YqMbmYLdPQEPD9dAO3ZVCoIeXCCSZZ
BSnYBj3h1Yz2Eiyqd+xGU88by0Ir2CS7g2aXwG1nWpmcEuy07l9CdUYx2lYnKNNd3fpxNpD6
1ICgAnrtWUUCH2rCrS34TJ1xvJJjvnilBqLcZaelCbM311q3bA780es+BMn8dgQuUe3iLYGx
V/Wjdwp2xxBYRazIPnUfeDTWQErQu9YLyLuBJDzyZ1hmTf4abGeMaheOXnGyyiOHjtfP8kmd
rnK1V0irtppviQsyHuwtc906q6Jm3Wy3AC+1NU0in48G4Dc0XxsJsD2kvJSCpsPQc71rcDDg
R9RUwXtykSZ0gQWpU0SA+h23TKdW/n7WUnwYe/qwH/uf/nI4tpAju4CACN8gmnqYwtMGfvQG
eNVo+5bLOvY1gyOvMPBF6qQ0gIt9VZrIBAq+ZoNm7SzfcuYWHa1Mp2mvNYCof6i46N3o5JX8
IpCb8geoh5d3LjerNHFYuhPL2+WZBAw5bICeiDY/EZX7M19KTenQCHa4csXXidsJm+gnnv9x
eScNggpW5WpC8MZ/yfqbc3JIcLgxoDM5euJBOuC7FpfMJOC1JkR6KQupFBdFA4MhcCMB86UN
58j6UsGDDi0tjvuxrIV5hsy/GEqeYkA0z1AzWt7WmlZ0w8phnvjHcHIm+SDV6sdfmIsT2/pY
7sMlfR4WqXf8xjtLf0BGqkrAj8Xm5VRmdzK2Z1asOsRdOcOfn9IrKqnIhLCC2fpMpmFnFD8Z
fDOpjnKLPuUJM9IlGSu5EQlET6ycCx+XZ4Tj98LEupnfHxhlNWN/Sq9Uxhj82x6HUbyb7mJH
Ymo32Nxey5qDSROPLI25ba/jh2oGzHqQu17rjlNx2v7uhxe7V6lhEcuB2YGkYHCex68IXKQo
Ze56qjMNs7yosrV4tICMk8lLCD1MkeeXnrRrVO5Y9wWL8B6pKPcvdvs9oigPT78s/migyRj/
Omg8IoIkADhinNQ0W1mTJPkJPeB+tjpIjEyuGNw36fB5x954DlEGClbhcTViPnAGaQieQUVd
YTS8GvE+iKpenrAL8xCA+RlZDyIs9afnGHAfx3eJ0hLa8EZxVn2dQhc62eR49pK2c4Kya00b
tK6suDxMsTn9lQ7evPzPR8yYXUnE8f/TB6YEt2MmWT/H3TTlSJU3lKXoZzBd42PnKgZrl8ih
M6WKfdk9eKx+sE+FR3gLOWjso33gh5YL6n2b5xSOrVXEb8Zb844T5ihILyAPsIjJwh6f8hCR
Zbuf3/7DntTCGxmTBbrOfLunb681wT1bEOZh083G4GRby2wBvB/LUHzERYzL+wRGj+DbnCO2
pmLepmC9EknK19+X6InfU0dhwtL3c7RT6UKOKNVDxM9N7co4PMfGk9H38r+ZBtA2SQKmJWAW
eO7j7D38rg43zC07kXSeRBo7i9UK4QLzPYMIj5XUS3zKuR+mZifNsTK2aEX+rP2EFmwLG0R6
GCLdM1DV991Q6MJSfpZYmvK0IyHYAyf3VVvy2nt0rW14XO7/8AxkSOOmsVqxLJaOSfhF/fpy
yVtqeznty1PP7qLgx0hy6BgeHYgF84uc1tLtKYgaH9NtpLaEH6g86aXcnUsn0Lw1mPk53aB5
T0TNii2Gr2N4F24WRkh+8XQs48Nd+HvZEo7j+lURkvUcGuZ5k7ghM+qQHvrGSZ1Z7RDhRe1x
o4NUg0Oef5hPK7WBa+NXyerzaygKiqKOHzMxei8r4xi19Lad+zmrC/2D6gpGsEkx7eohiUJ/
YAxvKw2sLN3/YmSUbGkPwfHeTdhYkW8lZp1iYdKSkO3n3zfyraWVQAfiQe9/c51iKbFPd9Bv
JMmZch+fa8SU9DRDfwXPOqG3wSj3ecn/YL9Cremw1iCFwEwSFSghsvtqXyP84+EmL0OT0jMz
4p2cE6kir/hhgFmAIqztovnBTxm/fWZM0BdTCdSOSLRsuqSIJmTPzHTADdsR/Ab0cgzXG59t
0CwcfW42g6M2TVna929pLQQz3fe7wErsvB8g5rgzn0qGZvlz1gbSyHpjLeYpd+uHgYKhJaYj
nsD3ophVlIT3eiNCqByj7uNTYHK/VWlHCxBn+D1gy9d4c+r0p0D29pgN+ksGNwt2bIEaXkLp
8c2VfZYIyETNTbc26OJpcTDSt+pibgG2lLWym67XvawSgvyYFWbMBgBvuipuoWtberrqixFQ
3KZ70tVB5wlAR2wa4QbhdV1Zui5PwJ0nA0Mm5Q8ytZLqEkap6DuVPsYjx72wdck9ar4h675L
dPt5zKAl9PjF40gI/w/TdNkD0xAarq1gHSr7HguS9blrJ8Ggb99UvisGV32WJypEEQ7BLzaT
uMzFsxtH1plRQ8+GvBfrhv6R/pWkEf3gNWQZulI9zfdAvu0cVj5Nac0y9QeG9XKVmGaTM2P/
DBv8kH1Viv2QrG7svca7rrYrjExsGHBPhlcbYbMhNqpLp14kecehsOOWCdp5+gCACG0LUQ1R
MJ59wzwi/1bZ0+dKF8ap0SRRMg93SN8CpESlz1wMZmE5OOZ8GV89P7vsXDIdBc0I4B0P1Lg4
FCfyQpDJaAnYOZ3GwynGtCD+o+tjUrs8M6aK7G3I7pg2s31+kZ7Id62XA/vXgLlg3s37p//P
lNtKn9NhdjKROEpULz73lz1l+Az2glcgcWQMme1PYTsbS1jsUjifdvmsHSj6JVoOv8U2CRJb
CCkugdSxUG5QPWlE19djyb4tCIVP5Bw4Tz641+B+CLAX3dx7CrAexhfERiiZPcsPDAmeHAbG
9kII5PoEBf3nPHXviqsJxGWOoutiMcLF4zWKxOI83k1N8DsvHeYi3P4MYrUC3tjuffye29h6
Tm3bMdJfXG7NDtrdWePRsbfGq9k/D3827fHRehMcmJwk4RPsaSHIPi0VvdvbX4486rsepuJ2
ZZGnSbA9YZ6B4fYxrR0cGGPXEHiCW5LjZQHnvgFrz8tSP8QUsPGHwSu18r7tzWH9VmoYvXl0
unIO4qgacM8vFADMYIVxJStOLYeMP0QAj52wfK9vPD/W7WRFI2qt11WnqLx8LGnEe9c80lNm
uBJbs2Ui2NDpA5B/hLrEQck5lsvaoYwfTM9m/LRhhQcd04iTvtdCaMo05u66nyhPsCi2d1lQ
25OOto9cmdVzKoKPYUAebY1LpHi3NcrtMiWSIX9KuaCKG/m5p+QccL4A6j1nTt6dZCTIm8VJ
Td0I4VLX8uomQTjybRYUk89qNlDrgyZN50yCXzDtOo4ublOSclse0kCTBOAE7VEd23gRrjxH
XdQ6FwDajw1VW4A5Ypim88pyk+WSoyYbCrnhki0+tbm0hobOGojfmSITxlFD27QQowrKep4b
ljUTWA7F78fEq9Jz/KVB+NckRPJupgg2z/ggeT8wP9CdTu3457FUwxmuFDwwc4iTDERKb8lh
nEWSbnEW5DmcO4SJMraQb9FAo88ka5zqMfniDzamKcm7fSEvNoaaWfc61i4SWRPutBWuynAl
IQAw1jlK+/zQnrSAvzEgCtUYacGtIYQKw8Qhio64wxIscjISZBVm+7uP0OJffDCfR1MsqFUJ
ILvEGd3H8kW+YfGq5mn7AqBeoUL8VpS3FzN4Ffp/DvqFgx/sOAMf5yYMoHUXqX6QKmLFRAYM
jT1T0WkLQ7jT1b8h291GF0zm6WQzmSOHK9X+DW/5w3D4wbtgM8XxUQu/s1MAySUa9frZu8Gr
FUy8fyH6e9AtgsV+pZBuSyoSAsfDnechf2OGt6yMYYtAVoR8E6RnmeMYHSbAto0lHWOEpStQ
7QvnH1mZAgUHezCWg65wNy05cZghM3i7gvfo3fNp0BBloGO1vnjAjzzOYyeazYpKMpNWjwRW
Hfq/cLcuO25FqU5qhmtvmiGXrFIsgUHGWPcMr42i+pHHr054owz6Lnnp8Q4wdTlhO08BxCFJ
fyq89XlVFmXZEGuvStWZXJjLxtJlDYMVFwRuCuLrf5fCKcj0waWspVsChx0E+d5ge0QLJ2z5
atGtyZ1J9ZB2cLnJfYfKAe+I3Sj8TsZoxNkkCLFwaINvNv0Znz/3oJOiJcmADTqoxEAzFZ9q
koRZP3+BQFAVgdOArMkB95P4GFwzpmlOYd2wF7+u+9cQOO+7haqwUvxURI3BgW0bpkOXqIny
fWwLhTxebFy3PzkDkEjXopeNpU2mHUdoZMFCZWyM/e/GgLAUZmn9kFUmGRYvizPQdLDOLXrg
o8MeMSjPBIuK6n8xGAac9edDEPJjZsVSod0sodoP9/8hkCJHInddPocMhqMfGqETOsLIvVnh
m4eXHZeogo6A4lfdCOUe4SbGUUYoVoXZyT0wNTE8vIiFcGxqbZ5XvFijzHF3btO9gBbdtvaW
WrdWFp/CX7nbU8x15QdNgYyNeHINboF+yGtpBBO7+ng7BxNoPD8ROhL5cLmwDqykX/iA3lKa
4RlBvFLiAdY+PKOvvZNWyRFaJ+M4X3G0rzb4jsiXqjTuWdSBRe80DO0kOB/2jKtO1735dSU9
QNgNWcdyQO7RpVcyAB7dMU+FYaF029CwNbRczxrxNYRa7X8qO0i607rlduLqKuIoQxC0JfcU
VIhG27gsFnayOTz3N1MqQEOaZMfL03C0kAsomBW/HqVO799BhUQSlvB/A5sgYZ2w0ie4G4Qi
ZE59pU/zC2Z0vmy2b7S/8YU5FoDTzKmiZXvQrUQTl7ufhSvP3QojibRuCTC4XpG5I4C3B1zb
7aKxHcjYpOSElcf8cGHf3V4LzjOlzxAWPdCoIjOAQeEg0YxBNvNYLLI/IFXpHYbYxWIg1OtF
IfgsAjk5iHMAi9cE13/xrSFnhFSeasVdkEDJVjNJ3YS38qHK6kdNyEDSDnr6U20SoytyRwup
BfSA26WMviuPjqHV7W6SK/ZpnnfBFxP/1KpOJhBRvMAbp/7Zlb/NGzK/6xuFEi7/1XmuuEiJ
3tgzGY4M6HY42QRPFtSohlHzzV06tHP0xgWXFhwxV6oQCk1mtmcv0AN3zPDHiJ3YvZ+by0gc
wYHJOWfgnd6n54nvg3lhJOc2TrkuqtiZ6Pk94yz832xL9Cw0SEdnacZ6LoqGUKvvNKBUhdWZ
Req9UPgJmda6J7KJciUStQBjo4Ul3HaoLbzAWohwTAfO+BVT8Om0RlDyscIsxEEWsueLGgvv
G5jMfpBL9RZ7YzbtyCh4iacHzSty1cjDscNJR7m3u5HYPcBjBytPStmW3EUz/lvt5JFLb2IF
bfjKgErnUJGNfZVXIexfSSHoCau0djQpM93PRw2sQ8buOmUqZivI5sMwZbSRP6nvg/27v5mf
gubD0mGB1ONXqkCWq4Ma6wQMtupl7QLqC9dX98b08Q3a3KVjcMO9Fw0CBdEa7GGmyOJX5OoF
zwYonjkb3ay/+ore7wBqs5AbH80d0moPO7OIBVg8p++2oigSllFDpc3oTl5rp4qyXXeypC23
MEZAj/7vk6DuPk7YU3z0eVfvP0CNCJDGjktOraUodu6z/SWYThPlgPU4Qg0Hs4kU03VtYAJt
NXmRHNuhfMxVuavwRsMYmN1f+ZL/FTV6vKdxbYAscj93uxWsfVitV1uNr1r/Ypa6nkLFIfKG
CFnicecwZAB8zuggaqyvmncDtfiaWZbUhrk2eln67q21Lny1ygBvKsVUwZixnAxDYRQWtoEj
7MHbVTX6OXBH3LaS+3fRuOlPOQOh6t/Pp0Nr7OJYJCerT9JdfYdqEOkPveaks4PAScU82Nzh
ifu+XSK5kRVmhpxCkagQUyyAlEqWMnot7C1dSBQA53sIFrhxv6Zg/lBOiVntlZ7PCkqE0PGZ
zOpgudm4sjX3lNlfuZvXbUg4Kz3FNJSQZyBUQWwrm3rHMLeGiPw4tUb583ee9KTHyxi3t8bQ
L0plJ/1sn2z9gB6IVjP1LqAu+XfwFGBqFWl3XgkC23C5A8JJl9oQyEveO6fpCu083OkSC1dZ
xhM9UOqi2u+WKPB5UzOzP+9Y129ymHVYxIpWk3m3lwoIhslZke2YGaDOPYh+/LvjvGnrK85+
kK1W5f781FvvxaluESnrcrnQ8gnfp0SzMP9JxxwccBFKP7+Tki8JHGgYsNsh0aTnajpridEV
NLyHhbsKDpRASYDnug/E2evWLDXLhwVRxRzUGifR3JcQ1MBBBdttq2hwtYw9E3dxG6Js/vKl
ZFxvfo5vy80kfP1Kp6mtGI3Mu5asQrpc1Ht73D3KSe9pBrz80dBAvwxcpRrjQskCBsbypTQp
eMXYPDrgtGzMrBDZF3yrPf8z0R39eEZwi9e5IfAP1b4XD3UUpwsx6+vzaeku77wNeS8KkrYl
XTu66+ze7Wwt6AvuPPsAXMVQDw24tKAsZ/8R2NOWnC6sb4t0F81YSzwIDmzVRxpmelf0IEZ3
voW2luR5uv6kP6RCzESxKdGeEiv+L0dfRGAfpqtnytLzmvFhEbIfsKPvIeCizsSqH75XBVWq
GDise16Nwh3rgSL9KSeupZBE6UaX8YP4UwNi5R9Fmim3EatQYU4u4ULHDavb8+IXwwh5RGjq
cfLREZzFLbAmtGTuLnZ0gX7dWF1hs8NtMRdXRujjS2np0tWrNvuqWKLudLTMxcIUrbj1k8H+
abAeJKKze71RSJYKfmbyjigJwC+4ch9wr3zu1tB6Akf5/n+8sYDDCO4BUZbLC6wu4CzyntDY
7cp+Rbjxn8UOk7y5f7J2yixkpbG9TwMlLXH7sl/0fEmg/0uicVLpn3VbibLGeNKSdYo4HBlU
1dGfRj3UF/b6MGDwaRpK2daYnZJTHt9a4rwnFHo+bNJM8wjx+4dVMMFT9ZavKp7mtndniLn6
u09fz+EZLOkn3TRx1vK9/qxsWhj135y2rrI8lmiKpJlOPjblQOIyMJqPJXvVtaoXocwRdwQw
790Xon69WlpQYLzxNTVD9Q/UNoiE/E6N7y4Mri6hHLiJpKv430EuB60mGLiNu/MC+9FzXTyy
NWcYnqej5lbkYgjDgunC6I38c5GJVt8XhWQzC1Y6kqWzKKuFkK0WPKJAnQlh2Uwk36D8znII
T5WCdnBJ1kYt+VuoZYDj2by0vry5kpebB+7vTyyS82bZI0sriKaTV46Sm2ZJfa9xcCa8q5j+
34R7iTZP+n6eASSZDob4ujAOznZyUR7O1mvso5i4HOe8JbGbmsg+ruarEIMC/hlV19cCexj6
T49QkJnjaRnS5Swj65fcvRgOQfJXp/Cpu/PSnfV6xjz7MCqQPhvpdpeI97kosez57+UzwMwb
H6Vpq1lVYoKmh2VivoP9E4ZYXgcd5uYx3DfNmH0NriHt825X4WZXBe6Xo/utHrWQwDE0HQjP
OvyuB8XpHECRXebcV3BpZNFCwF3WepjMj9+t+1tYzv/HArv4Cl/uXOWFKrFWfpgoIUd+1dJN
SIfr5IIXdMnF5Co4d3+kyi3RkjBsNA+2FVSqBPfgUW0TJNp0AwKJiDXdbO4pym3KL4yf9YQr
MMEVl+fQtrvQvApL2u/6Lk29O2H38cpf5I5iWVGozOmH5pI1C+/CeDZtNIdukhoajrfI/4Zy
geyLRKCCMJJMz1gMQXJUjkIh25m9APxYLKIGcFhaBXA2hm6CgwSZ2ni5dB4rDDxL13RBYrk2
OgltT+CKMAjYiOExMY8xFBW1wsJ5PhQtCWbhbtIbTRdWE+Snb2dAU6Jrc79z0fghfBRImGyb
0bfjOv/Cjb+MZlWkDSHbVoFYtphfFhiNQh2+DMOKq1wLvKK99+rDYfU8P32HzpXyYGR4uK9u
5PmzbvyQu/ATp6Ofvc5rN6aFh/yciZrglcKt43UuI20cFqFcOLyj1WN0UxBMVUP792frIGOQ
vMCSU9dKR1R8EO5nR6j6K3wShBuIaeOZohbCyqeAPU6Pb0G46IscDtq/ShccxdNLYwbJJavb
GzpyF7HaAolE5Znb0Xej8iQYrkhiJQLoUrD57g/4SMO8l8bafukALIDwghDxrzTuvUwPhwDi
PpJfyswzzzytGO8qZuQlZdpPeFfTdsXrdpl+bK2j1YzHlUK5r88ZGeABAphwoYhW6pDM7GfU
f9t1G7nBraAUXco9x9FP6E+HL1oRad7q9YaZ02XVbB8LWR11TJeizS+TjFQmJEeJorQO6mBf
tAS2jl6ktAZhr0qmdIHN21SOfvjSnOZPnuBukH8hN2SqiOWQM3V01FPfB1BNTVqpgBWY/82F
RRXQrydrntxUOBPOo3RiSBubos82K/+FwKROt2ncHs6aHPlxIZqTwQAjRAhrgY44GayEORvs
2p8eBRHoUmf6o41aqciOXieQYCjCfX0Z4flPKK6wO7wBadSldhkIq5iLK6/riq42Afi9cly0
bwo4bMeeC4EJRFXHk8MK/Cn3mAg2yu4jJ3RGEywh72pI2m5E0CdqVk8VszQIjyoIAInjUMwX
+xZDoVJcd1xD+If7tEmfhiKn5NZM8a/N/Y+TifAZRGH07ghf3Sy/3/UiAr2KXj886wDlYVkG
X868sE5Ot2ZYQ6kDVQcRsVo67lEfIQ7ABRSF2NG8Hw7GMn4ZLfz3jvB8Zdf8o9Is+M8i8Kdf
6bVRIwGiTCzfjTOjM6OENzqmbJzygO9vEvZdeVf+8w5rA/M84zCg8WZ5LynYdPvK7nVkxT+B
xDKjQ39hzdqg7T5zryr0BfqiYQc8ZQFTcXbsiCfCO2KnvywLZf0HS80rtUkjCZ4PsvTfq6+q
xezqxhAy4OIB+2fLU1r1uObANLarOc2oQtjrtzPMCLVXtSqvgbPc4u4VvxgklyCvtHNSJ5lw
RRpK0pdiTSuQ7ZBgkfwOo9oJttXZyuPj07tqCMC3NGLNJ/ZJuyHUV/wz7/z2/uf4p+x7Fggt
O8kd8WwmsAYNS56AyRdD/s78HArdXGgdgbwC3WJE3Mmajy3Fywi2JM5xj0IpfK7mLsRSW5QY
/IBElmY+HcwaID54WQ52b+YcSL6MCrGYKqNSprdeIcBf7K7a3RQwsxOZZ2uiowAl9BsCw2Vk
GXyAy6Emw67ODDULDCtrBk3ve30Z2NeUYon33c607rP3lQb2Ji6zceTOZYm9WCLB44B4HtM3
0q9AJUQTWaAoSMOu3hXKVOI5OkGKmGkwf/UTgGySRfO1sAZ0h1penVp3f2WEwvTnYY2LktFs
/KwT6xW4+jryI1wZ9/EtoErPZXCu4jcyUlMQl6mu9O2b7svWBUpnvuHJ5dD+nVXXyqVE3JOj
D/p0CXpC8DztS0M9vMGXzE4qHU/qixnBPVlXx8R7ohNFel8qoerEI9+Ne0eQb7WeCcIOoJ6o
yovip7WOA7OHYDjSs+gTYlgEQKVTp47+Fmzr/+nkE1C7isVHEO8W1Ns1jou7TEHJOiDRR7cW
zZlg/r46FyR9Do6arup8BF8/1/TGSjn46jerFJuidZ1ZqQhxGdketULvh+/0jB2UqMPcuTh4
oie6vCcx6jN9iSSzEfbGWw/w5yBp0ExgH2stVY0n//o2Y+ymbxE1mQSAgz+L2qp9a+apRH5p
VpfT4sv/6ryTWEH6Pt4SMgvuhtkbCANm59XJx6fgd4eFq0SgAgdRHXQ7gPV05Y1h3LaAUpZk
brkoOh8lhyueDzrwEhiJSxslVRV+WQM6GmL/4vnGLgZFMuRmYLEOy/R+Xw/7KTFrmiCoEWqO
h8xUJQftRiiFLR70Mr63OtO7mjOoHn4LlHNKreEl3/9QgPSTIIr8GDr1RUFkaOGE6O/akQvv
VLQE+eR98QK4NyEDbl7nrIVR1+D/n/NuHggUgJr66iQwAH71U3moNHqu2w7FdAlOrZvsrNmv
E0f8RcMdJOZoXBC4Fp4+LbXP3nbzrusXw3Lpw9RcIziM2D4gvyG1Z0LXZaMou7icwbPhBWh8
DETE14J58OtGB45EA4RiV8mHzlnDsqi/xpOviGkgqmBIRzJc/CAbuwDL/IckqDRXHj2N9ySf
bah0zfw49jqSz9NSwpP2wTxnn6BTt/cfuZeb/19TVLf+mrI5wpAynUIfC3mJSnuAxjBLr5FW
CNiv/t9LtK99dJaw1DMSQknHoorBZiMuyQQGT8lo8JEf9cEFOXTxw9nxeQXibDikG/pds7lZ
GBChuLwjymqm+ZuA8dv3ZqP84jm9xeiw3GHuzsUIlOIDzrydQvMbUjK1oLOJTZZtXk+qwhjr
zHo3Z8cengboMnY+wVu6v8TQDbi+6vKB08h9ALo+mLKtLNzIVtslzLtwuebDvq6v+RvbiL9a
2asQ+aEdovr8+raPZuOO1CpedOCzB7TEMxVwL0pmtmuiV7LNOV6ll+AKhCGgKtaPIWAPp63R
l9rXhB7KN2vAwUrrrFsaFPxNEjcXazZW229kAe3k9wfsG5I0kU/6dkXR9S0l3F96/essSqtg
YX52P3adlWu2o4CvGtbJ6xexpVhiXrjGyZJLgLV+SxsNUklSjjHoBrqshoSHnmZMjpVCMP8m
DthaNcdJiMZPt+YgtHFpsVvc5/HkdI7nIwuraj4ba2afdkTMbKbUCNzNNikDwrE+kBKQEo4w
GHFO5+B1xLi7KPwkS4JnDWSwjHln8l6rkOap2a0yLAbJvXTXp6m7sXyNAAJphnP7/opKCNoG
EBksT8dXx1RMQ5U4OGp9Bt4ZQ1o7xZcOzaSdxCjBlF88qBldnfIAviN+6k3SVYHZz9lpKZQs
bkEFfR+x9H1wS0UZ6DY+J7GMIFOt4Njstif46zSJ3XhjOrETe59csvHlYGdf7F+C95ctHWHf
IyaBoRh7bP8js5fwN3q7wY6todMoiZc+xSoNbHbGYiYNPPSkOrr2kG10liaClAoIv1/nK2EQ
K4TdpoQt8DZAYWw6qhgo81IQl8opVHDLjnwhw/ncJAQuHSOPOROZ+z0uTdAIyej28wCP636F
KhCpaoHxQ2R8j6dBSUKVzKbXrjuO5ObdrsyWoGDgHYCFWmHOhEYuWoZ9rlgHk73soBsff5Oo
XH+DHuho7cZgLF/YyJL16RjCOcaxICAbpkQnQmOS4TPdyTYLiuWMiiCs7SyNDmj0qClR35fr
chx6fnXnwIL5rKbkL+FZcexz0s1TCck4KgAPmnBwN08zZ0VJo4KukNoWZwnQ6UVIM5G49qIU
JOq2gQI7uaf0LJ9UVZPKn59eRr2vqUP4NvMOz972tWxrwY645TGlyxAaa8BYwvamlLfCo8lW
aTqmt8tIX5dIt8duun+u/1XL129n7U2eIS5BtaKLjWYVJyyDYvDggO19yaydcRBFl6c5b4aM
K5l67F3K1MQDIa4v4SVHwBRmOe+zFaNybcOcDENYI18piDVxESYdaDtuTddY9/6n1XwiJziT
b57WfDlWNggtUZ9OBdlfsitrY5/A9nXJkrICJM5xciVmBe25923zuu9vmAyoRhXYd7Gt6/QN
lxZTDN2iIlNjtbld9C2qTjHMGQOE0sza9mKNA1swYVzgyu/1kzPSIaoHVya+vLHrK8VIsOCA
QAem/WTtbiVkEA1DGg1ReLeYJyOEhKVpQGUlCvDfIkwMNAh9ITWIzOWLwt9/gCOYUx3s6SCC
JWVBwLuMOh+DhNAFz5wTcG0RTgRmnHs6BVJDadEm4m+R9DPhLdBhi8ftuZEmnheh+R/4/ww3
PbOwIdRB4wlKU+xFmpy41WIXf5HmBU2ANRttzyX5qg1taljyy51LPRFLeTtxSJ/1IiuPyr6X
g/DHVosvMQxF3sA5cYMQ+GdeyViiHbTm4budDUGMMlHNea+MnqhDRcAqSdqkFNo8yNyv/AYJ
xe2YvTXMpCQA4uLHJytZlUiUFajIbGOaUtzRRRtEH4nE0a7l6s95zPYIDTPSAA3OdNwhNHbD
2xY533D5uyjrOEXkw5qSxOLMyNyBHK4ZKJmqdOtxyFfUKy6KLvRod8b6990U8JKAonlt12fo
6teegKHSox9I6wjITJ7dqjN+wSL8tpHM50ALmCeXb2BmLAugl8Hs17kCeZpnVgCpE1wVRuBD
QFhwAG3MVPLijJ13JNhcTYBAuFUN4DITpBR3mFdjp3EJ+lmU7xu22fUMgYDWyN7egKKz51FW
bBvXqHEgNjFGpuoa3tGE0Y1NY33D4nzSA6vfg4n/+1Iyb4vrUjbXhPeiWWeqYvpi0RVd2XKW
gIX7hCv/4XkYWDD0XVXEFViLLC2cUetcc3ryURu7SYNpfm80QYF5sB7kaWr9clCjRrqcW/yU
jem9oWTrT2xX4tIWXwcFRl4DJIvTm+GBb1F5MMjfoxy/lshblKfSHQ/5MpovOKBGposbLQXg
LgBFoeOHAwIVlVLcdHnOsHoIk8Py2fSfmqEQLzBRgHB96d3TrkKXcM5xakdd2dUHzVkurG0q
CJrfRV85jC8ynSqB/InZ3jGL8iUfLAC+WtZTYtCdpD9ZktI1HFf6vuQCSC2vkA7NgMeEw0ek
HHVXoc/3jMIh/gtmznK6MHlKFM1KBxSoqTfPQWenfgODgu3d4jA3JhDcgfPVCeBfQsoYpevK
FuSMbNCjtTLGlnGq5R5q9dKCfz159NMGI5fRecaNHF3jX+A/a2Dmt1WQbWnHgUJgZjrPQrtD
SSf3abRGRqoC3JCb54IQOU9q23sUf/lZKwsn+0i23d/xeCAAMZaNVBAPGD5dCYhRxOAM2Y/G
1pHXyayfwa3QrnoydcB7mT0nWFA8NtRBovCqByNOhtRzkynEpHa27PwA5PQstwIqMCi9j+CN
hvZF/fPfzrGcx9estq0FgiIS6OqyHg2X5KIu4A+XvIBcDcZDFoLh39Dy5LOWd9oot46GBrHi
dJvCQOPoP8+5wf1p9bFxuSWA+YTagk2fWom5nlwXuQT6udibKP0XSKhI9un4ji+o1IBLO14P
BKaxRls4o/NzN73u6z0WBRPP6/LIHdSejMdOkQKUezGQq8uQVOA24psT0+21WBL5+AgwvxHP
NS+g3/QaBgp1FuVlfDiKDG1wlG06Jr9a+6wF147toSbYYSPZTeWfl/Rd7BaKjPd3ZdVmC+1s
LFbjO/a8jpvMjkGUqUSUACM3Di+oFWTfA1yn8IEq8ngNoR2ldc9Tj8QFNkg4Et4vFr5FpfTx
p9FU9R2iFU0wXYU9PmbAk37pZVu3LIu6g16J847EDw+z534aUD/k9duXzb/alPm0TIi+Ltvi
67YwQhPGadCBud5gDgA41ClRp8u8Zf0rd2FXAZCNGgZqInw2oFlfh+qMy9lgiCRYbf8gQ28S
PkM6n0zMdiphy3bGeyJPuIL9kZOUSgxWneVS3p6eyC+grL3K6rwATS96uONwlsztNczUyvCJ
APJiS+/CnyQoYVNjvIZLtECkPorN7XKWebD9wm630XPZTCL8XVDvgrGk1uA0MSDRzGCyB6ND
8FZ4hTgDfZobaexxOktHnRgpWMZE2cm6otKvPvaxgIZ1oYfU4U1DX0rPILLg0LqQLdA3Ik5x
OpwNEN3DBBmwUiyGXtd4yik95aajY/qMiSYFxAbSCoJWG/NNr/dv7G/HS+2N5g8M6Rmm9mey
1ozm/1oWpDi7bcRX8cKJP+rTT4AZxORbjdmu4SwNN5VsU6mYx130sW3nbNJbXYuet2lzMpoB
LXPqGYQPEA7a+mbf0C9SR8GlAdlEmT3Y122mA5oUjbAIlIlmY3sgrgX5/I7nkbobNVk2NeKk
HL7B/AYr91R8/F1h3gzye6Z0H5DF4UrFXWG2RIfVbKW2Ufdlf8d3AVWQb8Tnaf0NMgktNVhn
AzR4ak5nXBadij6L2MYH+UNiEX1tSnVZFkrnWBTpi/CC6MMlRaxrusbOm5WOVX+wXIyW6NdR
MqkN1sKBixHoimwkTBcQdpjje2QPByrtpD9MX8VIxIgPPL4ahd3Yt2CsQVErHC31zFjX9S/1
EyfXuchexU+n/3Piyf0nFXSB/GChJf+uPAZnSDcU4r3EgUrWJmDxteizDBKTljKvn+sjPPmV
L5n0lyelr/gyjoX6GVVuvf5ACvo+y/8zk2LOg7lkfgXs5EdZwqnb+RoEqTtsK1sVupm5mPmZ
t1gN90giEu1mWghgUfDxwVR0a+vLSEfS5pucKaPJqSInvgiF/cEgC2hWGcrgqo47k8xiAlvp
zEtf8dDv8BNOdtlY0yzEW28KVVwBfwb+5nE5ZR3V7ssX4KbHk8q9hH6gaA3gfG1AmD0+b0Vp
FoUN6qNCi+H9utwpUDknWHtP8hpbUcFdN/hdoi10XowayhsvUh8ctA90bwGxksnbEjUzJyTP
M2+St2s1RIR0SFEAkfzAtCdNueFtX1vyS7llLkzIDKQaY3xc3qklFGuKF9t/tgwE7H6xEaLV
zrKzHhA7lIg07ZVrxkdTwDQzXS8X9xaebShgGp1aYTKfDi2i4TMm6a/ME8+fGWYvOQ2FhChG
A3K/4CtonOdRvXi2C2B2T2TjPoLuRCd1fzz24HCQzkG1iZtjND8njKzmXV+gcsekBsI8SgU2
TPMwrnJIybUaOkWKFIeAigtxwcFXXbQFCECv4MDVzdgNCKBlnSOzhvsRUq1U66MyHkM1E2n0
NCj2P0gbFS7BP9eG/Qph3K1t4nUazvDPbglYO86UETtL76FcV+THw+FnCjOiYHhLbtvAbNVJ
pbTN3xY5/8BDoWyOXMrRf07HpOQfkOdhwbGx2vTWGRtsL82ihLrTa7BmkWXemtZ5pmckR+h6
CBjzbv7x29uFJrWD9A/VwnK7d6x7h8t1aDEfDy++ZpGI0ml5aBfhBC4ufY2QSojvdsc2Q2qU
asmKhGRb0SZl3bGYKEl+cnyD2ard1QgDmaXh0zmgLxnaThYcMtg49i1rfzrGqYunDo8o1CpS
NVhKgcNFYlKVOR8ruZPW04jI+ofw4U2xM8oxA1S9Cz2iTkmB4/JcpJxXInBb8kZJluQGJLuN
/Nqy8tujPEhBMACEY+r+rwKYDe5RHz0IxPT1KXd+Rc7QKT2ewuCPZrZSgpIl40EEROYhaK6z
+tFY0x6+nBu/v7PJq51dsDcHTyV3akIiGlVxM1bYOjaNFgPAgKkJmOZOC6kYRJCfoiCGJJwa
ZG5yK2LrmGFTJBmVdk+Umf+emZ1wqTeRqSMEQp97siRY0XvZmFqmXFeCtljwc5kFiuoKSp+T
T6EfBxhwAwy80f7+SGD4PMeynFDrBiftT9n70j14r7FExso2k93jIfmnyL/7z6Wb27GCrawk
KvnuYO6PK6YdqwH0EVklevHyzzRpHnuqzxAWITwWAACCRZ5tY6PakqpPvH2vcgd8x9onztcq
yJltmOMXaeaNuRCy2l4tAQ91yCstzAUzmRaXLc4eK72c4ROeZMN9EF21A5G4pf8P7XlshYb/
jFcJEpE8IQ6CBNDrG7zXTVws5cxeg7pvEKRtiR3rvJ+BXdZjROfleDYzzPfkqERopzkPTkNE
ES2YcLufabVM/HL1yCHg1rwIUjjPmfR/5Sxd7i06SmUiP8t2HiJhama06y8+vERQV0I7Zwgp
MWB9Oh71UAdzVdBvPQvrul0liq0yWYbakjU3gyx5W5FJusj6xCnpExwuqgGLjCrJJV5cXU7y
5qwoUeXdCcAbRQ3sab6yWf7YEiCXNS1H279P5r7nyyJo50UCt91BtmaDppHNbvMG7cm0xdrj
cB2VPg3lz0i10+oE8qt167viJLmyAkYBA/xcvs+JqTbtoO3yxA926+DYaBMy46RrUEHYqAkn
Od4PO3Rt4amZPrU5m0kYMR7ieMshe0kYG/5C0t7izFueCgue6yPyHQg9CgrNIb73xGMP7+jE
bRGC7zpcUV3JmhWVVdKLByFHfxLcyfTyKjQn2HQoweJyRhdcNayFoizFRsIjz6iD7wLBqy8I
YZHyCTSKStAL4SwrYRX7qZ3IaLrgMcSzl67FpL5JTo+AgG3h6/yIQvvf2OswX9LMF5P4vay2
sdQ9+yWiBZslHJuJNUc//qYwCJxZQ7u/QPciKX7depaszjpQsKLJLOdF2OHi/WcK/ABmeLyQ
mXu8qfPXyKt3zDNHM7uJ8Si+2mHpM/ad1VftdLMjJDs9ehl34KaUOhSlnhRuJ0RPI+3Vh6Jz
TrLBhosjh+tq74aCLVWCxx9EQOYwwuhJV124cH50iZjrhCIilbpqj9UZeRaHJIcw0bIdcPDd
ITy32ZuOn1vivHaz5nczVQAJxiktmdQKMhrAR6lC8rYSqLaSAfjZ76sN4ThR0mg1q+BPQkzw
fyRCOemcdEwuyLNKypLj101LQtUXNyA2aSgnR/7MXBqhIWp/vmfo6I+tuiplAFRxqd8zHEA8
fXOu5rUHyQ2lzQl8ZAYiwBov82Jnsod+yi1FJRvm45acP5ggkLT1F600q0JL8hvGyUqvpA8H
5vRnLOLFRZS9cnhbNIxzHzqh5TVEhBnMoVghibQ145PoUuOl6pqAWtZyESFGc+r/BM2raEG0
iCLuIU4NW6K0rAnM0u/HsjT61cgItvzTyhemaEZAXZLysEsJNqz4ce6EUiWZxJu/wkYOLx9f
LFUzPfGO1V5FEinvZ1uy4FPK0wFifGFof7pcVthrLQzOCTDw9Pd8Je5FbiY9cze6TQF4L4Ad
t1lGsbC+sTcr3rNK5T1rB4QTarUlqPirgcVLNOb2RrjKY25LiZ0RNqJhOWiq7mnezif2PDXe
nPDuYYPLh4j4XmBFLwOtpMXJ16wFXKnlIIG6Ad52xgq25XyhTtrnQHgF7fLCYq11EsDrhJh2
5aHrzCjoaQrvhKU674mCMSq0MeKSbKkMme6iCO0smHyctallUch+sXktUpcFa6rO1R/w+KEj
sCi8ySbR5Tq5TL1wpIyEgfWAPcvKHYsjX188jUqXDufSvE8sCp2J/GZrEkY/yl30YsuxdJwe
0xo844G8aSf6vRMclmlZLpub3QWG9b8I/fIKBrv5Y5BPvWNFI7PP5prPc/jSbcEgSSqF7gBj
CpC5HHPPmRmg/3GcygieAx9MlL4PJeFIvyy6q+qtOHWQtbfelOC57A1UpxOSY0nisCdcGLl+
cn92Ubf9vpLB7Aifb1e6fF895OLBRAcKCl/15dfq0cxSjMZsQhDuKM0p+A8LGU64QxEzyJfO
DuwDhMMNkluLH/UIFx3dR5B0vhIsEWARdK6LvqGaw301PPdtsJhHaBDbv3/flSlthr9e3jzc
HIfk3M4frCr5KHfnbMHkadmTvZcW9atpxxr3TUNwjUk22HykaBRsd52WrgYdrSbaGsCyn2gd
QBKArVlLVOLRRGl4Zb60FG7+PD0nXGjQI5gDkd3KsQxgWe/1REwXB2IvE7xnFBvOr6vwYKsf
2x6PU5X7XSoFgbM8pVukLDgUyUBmcFbM7CzKsTkWDMYZUETp5MRnIUhv27ujN8dsx8t3P/4Y
zByVmgnmToZQRAcqYDJZG63FBbMbOnmjCX6uuOlxt5zdzIqygqinIODnRV8tqwI/pBCAezQM
3jFAhTK/TnKr5A8vqFOzLYCxnP5AbJfzbrzXI3V4U7iomNcw1iz03K9BmO1jzXCiqgrmZ7Sz
DWu+7M9DmhFdniWevmgRdu9kCUruaVVxdSbt9FpXD8APYNdZBds8QnW6wERiYi3ki+mcsH2f
38t1Imeu4J57m4qNYmNGclvLEJ95oy0SJApqpTK+lM6q5abjGuHhWmvwfLqURGXCshBDu6Hg
1KNWhiH8TKZqlVtx6MwZV2Ub6QvyRxrxKjlI99RRSho+pAxQ8N2K3m23V2OnELMKDbDk2QpB
QbFZdQuMTyH360UinrgxN4JbKDRGzlIUKYbsSUDfvKz5AtYfkOZIyX4PFv2Y4TR7KnEvXbk9
U3HMx/a2e+51z+cD3CpcUUBAKlF2QqA6RGnNH2H/RbT2Q5Z2o5UE3oTQ2HgEW+9WFax87qsX
dO/ur5GTOmKZKlb9rWBbBIjJ9khZSTx2bjl4F9UjSwp+b4fwWzUruC5aogKEKHmKEEUMrRgF
bCgRA1AeYTKpGyTi5A5EXIMi3Q9zv7hPm/nszUUNmZLpKehXdfecjwy9QSjArWxsyPE+7mDk
No9sQGI2ETAYEJSP6bbUm7MMkFDryhtNxIMpMyDGFvG5Gx8WPvbpFmJ5bnqVKcWmzELwZqH3
QK7WCLKF4WyLSI2TCOHvghB9IwuaeSdD7bPtH5hbIDv8OcduPJ2iwyXVybjg7mjmW+XYd/ZA
0YD3LzALCPLuP9S/hZQG3/6Mlf6kq1cn03jzwUXjWfs0BlUqi2uDAE9CF3jw7hvieNSQr2lS
0K+ZbetAgK9TEzJgwrSeu6UVZOSqikgEe//C6kRwvozKMc6++ypoRM6wZGYYMKLQv9Cvg56O
5J94xPy1yqCgwcf5HBaouRFHf4nsaWy1uH/YpJ6Q/0+gjJGGMiimFw0pW59PFCodsJ+T3ToX
q4qWe7+R0+cyBtsiBwTM0wcf/08HDriaAnQgIMA/Y9YqVKK4igj2B2Bp926dqfPSkYJYKJcu
+MgJDqrIOhuPfVte07OhCJ04IkqsZ7cfsyhzuSfTs3nj9kaIzWa0Jao9icpThUQ6CVrPWWks
AOxkuwrAQEWlKAmV45NW8HI3PHPEeV/NpFDDvrGHIDMbfMyHiSTyIw8qT6NuuEpNezXcX6Q3
bqC5n2nk5CDFzOA8Liam022yOijY0c+sZVNY8dlnOZ/bxP12X03bSLVHp8dnV8O47fkrUykv
JVOSnN+LxXhwISqC09ZCTDkaEjQYVB3NQhddmTEQF21f/VDFWyL29BLBjHWb49Ht2WY40AwZ
aKwMoE7+3NDkaSQC8m8o+gItj8zVy7L0ir8Y35ch/jhVIAvweaQ5GQlsBKi9w3fWD6REPATi
ZseqFtCOPVz72e4nRQDaROJTm3d01O/zXW3RGEEFMN+LGH3l9e8CtG5qJfOHsgWVzfI3nu0n
dVj4+MvQutMJUUxAAFaW2+XtFLWcB3tWxj7wEv66pO/MLPEOjO5ZPOfLkbJPNkUyxNdG+bpL
JAs7+Ge0pK10ur+UFoy0qkmwqx96/uGuo06D5W4evzf0yPJCL4dWeYLS/Ts+q3TZ45WrvDM7
PBG/4zzbDIKhIjOrMkwXnSMgSEOn8vHCaVw2An+lF9hCQLm1VUMVBSgSzs1wmc6XZl+Opxph
D6yd7obwsqUDN5ZrDzw0kK6FoM8Z1mGGCa5GnNjWCUZQ1qAna01Mvn3lBlBUyLUX/qHaU7wc
XwtPl6ajTjlDCJB1+80ft14XJGl1hJXO+XZF34RexA02Rz77niMZyiIgqx2qaSvDMRfrdVrF
CafQa7F26G7g+7ZvCT/9bfsNPbsHABtkjULr30Xrj22iRzDQHr/L31AYR+MaKUCSdWM8bq0k
EVgiTtsQ6qba6+4LurpLtVWTlYln5htCwiqQB6MG7OxbQe/R7J5DzVYctCuqOOVXhc9X672S
iQK9g2xQDVr200pV2Fc915qP6RhEg8rhGoXHg3fNyCLaTUpMAVzgFCVn+gB96a+QHv5WNvlR
rFC3ugy/3ztxr+0uXZxLcfvr97kvz2LpsU22+OZ67QS065rCpgD1BW/KFwYZc+q1fmHm+j9N
ESwdPbz444+DdVOChqIUdwlU71+fi02DOyzQY91QJO9XAuAOhrtWwFkwGgW3V91i9vssNKHD
tMHAGDTU4AItPrM+zbg6gT75ektxPBAu/XbNmUAv7D1j/9d7yXMVy7Cpv6R2mUuJJ1+ZH9mj
XTJtmkdTtMOPNg/flg4CrZWWTUzWvwDujNI2T7/JTZMwvDe1zXxPFx2Q2uRnoRVS9laXVfs5
3TOPlgxo5ivrQViiUOwogEBxEYIGm6P7FPLnEBdm1qvbVIue5NgGTR5HBXorSPzdqHvMyCEr
SZ95+8r5E2102IuBzwV/Gucwk/2kS62bSy7hgyPPhdjL3c3ocmWxOEe8m9SKddQZx0wlioSq
qsyInfCMNPgyCRtc2Y5Uv97dDwa4KWI1rvQGrAg+JTqRxa+JTrctmm8KRzdMJN0WYxRVyQ38
3gtwApem3e2c7jlSnYD2Jd3QgsIbjflbC1ZwABbsXFWhWVDyqdfMPmKSOTBy8vwJ8qEvb9aK
qCgbRB0YFyD6NHK57kZFBezAt/RfeMaBGuv1cY58ffYhV8mh5M/8KlYHdJh+FtAS65oMocFD
0bMCTyhzsO696Yxvc0hp5XDbrl6JV/XtdFd+AKoWFhc0I+EPTNDKndYwipzSSx7tL9wdI8Kl
BGsWiRV2l3h0JH/dc7Hzra8DJ3yPXnIWotzPG3LgZvr8tLS+NClpi61+kKwu8lUW9qqgXZWD
uyZtqLddjF5isjKlHKN7h4b59gJVonnTPhqOXkG1hexj3iv8aS4QZJlsS2lileqivp91isS8
LBrr+LESEfyJqoqUDRcrXtaHfQvOH5XAfo6v7TaTqA0iiPKobELvPKwU0gl91yIwJhAdqPJe
iKkfZiZoLV5Y1yQnmRRggEuOxcEQYrA4njBxbX1yf0syDVcctS4Id3dMo6Hr5qGEp76kClZX
Qa5YzwTDsU48vffqGoDliiAIcASYIcV2MspRtxSMrI1odU2DXfQiR0vQ+7LisovP11TafExV
YsIchyDUtxWAcOuAeSWToQ3zsfE4u9B7c8bAIMD7EJ2l97Etgy0An5ML8pgin4NKMJzK8aJ2
60v7Vs+wmuesQVA02yvHplM+7qSqltEyrw7f4DeFWVfNsC6LlQHQB3mYSXBuwzfzVKMudUWK
gHKVVqXDwyw+xtUMpnwhtjwddT6uqfqIK14N3F4uG7Vck9OyQKgrntpRBJd9oU+hvyXGXt6w
9N4LnSGZvARGc6gzqVECIOwAYmV2DRQ0XQP+oRATikOKP7yoMbTsIEDktuHntMNlbQ+i0fAo
0HfVISd3Sbd3MjbCIo2UE6Rb+x3X+bLaaFDqtOxY5QQle/tmuFvSpVPbncafwVeeDR61Pq+W
pBDFWFm9Bj0BWQK3HiaAhSrnXnd57LRNDgfsn6925y/Y9fxNQTHkl/BLEN998NDwsmBedmDl
1Y9y7kl7rMx9F6n/BmoskM3xwZEF1Kxa3TnG2Qdx+63FSHgvF9/+CZa99m9y/MB+4m82HGPD
uzjIa0ZLUhQWtKMHqgYcS4lto3ywo3erfpniq08dw24lCbgGn0S5gxLa0NFtfOwwGCW+i22X
0kw6BP4nYmkECMDjAEzZSEepnDC4nT8I4uBwcu9mnB5t82BzQXtGQ7RKYr+W360Afk/kg1Ws
4RxIC8jQSOl9mUyAGyQh0k5R9594Tw6f8Mj3WJANTTZAPIciOX2MCqrq+AtP7HnjO1G+HCJG
aC5VNxLrcbL1zC/Y4DE4ykrA6CXpBtUHeVjLoyEVytDo56yDEz7gPtJifk1p0m2QS2nEvPRl
Nsvyue67uIbrs1yW60Fx/BP8o6OFf/R72s6OdRr36LjCWvk9ut+o8co9MuuCLaAaDgoHh6hZ
skIh1/lNNWs+/Ysb522o4Gc9JJWjZyDYfSyOislkdmm7xBxTTZd33oR0okqBpsdJOWqY7SJb
+W4m9zw1lPND/KHcZ2k2tM04H//PHDmYP4VZWrfsaId9Y6p6jCrWfyRgsSBJukdJNfFhLTlr
qJ5/XHi051vqO5x1Xb+wz2wycD7fEVXq9UWTuo8ACLQSMtcVBcuHbJA6iRbBG2DpstgDesfu
u6jfIKM0ytqFWtmkmcrh9jSJRTfmN4KjxxEmHVk0De4Fu9oaxRd9zwTa9SiCd56kXO3/Ir8j
JrYhypWbYnloz/Ni4wUg8B7XLQT4FVeHRi1NTCmTb5BofOLKQhpGKLwcNEVNxVGNO+s/qBMh
XqR5dR/BxaP9Wtp0NbzQgqzS9EIeM3v0EYNDQ2Cqv5VbeFhAidR2biggb1uQJof91nH/p7i+
piVgd+JNvrp7tAiO9QY7QmNQYXS2o/2N+e9uslQUG95+Nt4hiqXKR3oCU00/7cu4ir283OH2
JIzLMjarpj8rM4PAmSyaeJ32EZBhfhbqeO8ohW/Jry4nVS5kqc7CIoMTjUTcRKCe4Lqd2t2F
+zW5dpjs3P+lMsNzHPhZk9fTtZrqn2HiUh2jbbln+GyZiIVVX2ESBaRgyGyg94Bw0zLTKaIf
5t2rMX1+ZOw7SZp/EnIEIYtkzHdtD8MWuChZ5JnIlsmAbj8L3vgLNiB3v/9IWz0pttHBamUx
imZ7D4Q0599RUKMrtaRJiUSBxH89RG5K7Y4E4bHooSSr+KwwTf2IeaVofPU6jHuBVuuKgdOy
thou9QdTvogevY87zvzmyYGIuFylJ6D0jBEfYI23SFzP7mUGJTI7nPXj3l0neraUlK9xfndj
IJAXDbFf1x1fEne2k98KhivTT+ZoJy8ZO8lSFvkhM27+48tcvXvfpdqMNw5zVUrwLHaZHEA6
pstKsV8KFIuRxjZHMgFmJ27cKJXpNvs4DBQ8N83xo8hwGbMOyIR/MCaj7G6YBhw+n99AA4DB
Aq1gWRWy1bQvSoFBTCOOKvD9fqmqljsk4LTEqbx2U7sVJpeO3z9K1dvCN/8mQcqCn9WJEEUY
51MiZKy1olsGnVckdrH6Zr+i2cXz9y+CgZOgGtxA57MXr6G+sTH7EYQVVP9PRLgCcbSSqR3S
BamY3Jvi5DeE42PjdBjAspqkgE90UzlGITO6iV9eKtwtiOlgeRxCHQxqy2A/xHBzbLrfNztV
fBbBlB2i5fuxG8TKeyFizotPrZtwXkQklTAeQZz0MXwbB0reEFDpMu4AFJBd/Esps0/9YT+/
khARxG7EtavabS24W2cX/XENg93YfvO9PnxJLuJlu1duNldOYe7sm4LmYTfFOmQicXjfjpuL
FdJbNoGpStDe0sfX+EacyK1c04JCpua35Vb/keh/jkNTbMae3slo6nCwt8iohHcIETeqK4DO
drnHvn+sIpL6EXGhMzHA8/seUhMC35tKRhNKsvb/mehCFunGcGtwt//oV4TmzRSFh5jrklGs
vaULeXJJteca5zON/8h7JrOAT4vgDc5+bQgvQul1xHNY+n0GU2Oml1xRtjAzmBNAUaoLXmFC
3qW/ALQ6mWn1wZKR+WUQfsAe3DHZIHSiHiF+OgXn4qebF+FdgNmN7We4FKDCD8cePCqDSZa+
6KTtFle3+x2I/bnpcPrHirZkP0EfnAanLYIQYdjMtwnzQpoVuhLutUars7vTCkt2dB1WQTz5
Nnc1dOcLDJFgsNJg1PRkuZOu4rJJG7eIcfOhZhZOt3h2uP67rJOHo5rf2/2cfkPw0a73u98T
mQp4L2ymWxWkWmyJes+4xH+b+O8Lv2Io5MY7o+fG/PoW69UwdUTWKCZIQy7h/c+dJr9yLHXY
f0O/Sa4CV94U/+ZeZKB7RPLT4sSioya69VEZqJUe4B/bZP4FX+fkan3J4N4bPjWQxR0MipUk
+MBSk1WUKyYtL3JA4si75GbM3/LEm4lp7T8cIvPx20zsVAlUNa9Zu0atk+X9YIjQeN5TJjJG
HcZc/H4pKnwuWs19a7kYLJZnvGOXDzaPmd9NJhy38xQFjDGCP12fWsJIk0wF/LrxtYABsw6I
DbXg+KHN1E85h0/ie6DPEQ4E36mFxrm9SxNS8QZHUfzBQeCpQQrh+f+EEfek5Hl7S9a0IWjX
wUPp1nxa2lyiu4vrKLFg0t6Jb9FOgrHMHjLTzxmUgcYi5Nm9dnprjyzeEvzvqZAp92qCDohF
X3Xp4wW4SaUbUCYCQRa6WpLaQ2uD8cP282WFO2rOSE+6MLAJrvKsnwt/NMKwYRS1TAyaK0Cq
lbd7GtTcRx+YiS+Mticcbm8isVLsiBTQ1dIoNcCHxQQqeoJ/HNv9dDCgao6cRhEeaEbymOeZ
LMDHRed3inPBiqV9SmqlThsw0lTld1elIC8HR5dn5D+7nKoH+WzvoQCC+wJZy3O3xtMW0fJB
SRghotC84awHUn4RLrjgGvrJ7KH0ARzPVCSJgyOGX5z75gYfV4EJ+TMCggHsaszjg83+1OZh
vw/9DbwjKsBwj8kmYvudN+s1kw9OsweK4kVQ7JANPMYmEcV7/UzjVPH/Xct1cAwEhVYQCEhA
wdliUq+svPgLTFpq/V1R20FNstLOM3FjtjCzEl6V42WEhVwS95vuqoDk/+0nmTaHnOWuRuSB
hCICW5EPkE4SCJN7urwfSurTNfxVXIXFh1QYfXKXJxBDOrOrroSVli2rFeE9QffQgQC71aa9
pKUIcIzBc719fIykm5Qr89OP+XQuYEmb7qOSk2p1QPSJCV2OjFOQ2JQI3lY8rKVGhtdz39Kg
guUocqkJg4iYnCPYlYvs83A2LxdRCZGFHT6jwk54xE4e7QANWqByq+prwc7XNQEkO2oiC0bw
RdusnJGbvswgtR4FZJwZt16ugNt+8sWJ9b6sPCRJSZXZJZX4+nxqIM499MXAHHAJGM6TRSmf
UFJm5IALh2h+VEihqZ80B5lQnME7IikjnEfwYZQ5nb+ezsszPB5imn5f6Z1qWBEeQfmDneoT
875RTzZgDczo7t5eekYJ30SrpBZsRT+ZlLSXNSH21arzG2IrOI9Z5k7aznv8cWGePYBcQ1El
e2BpJQkbgYreJnotOcDc69VhiAU22Y9xxuCgg1vJ3w9a0qjkaj4gx3IRopZeSk34UNe5NuBS
anMVTODaAtnA0zXLIW1qQTNftQCW81lmTkCbF3YnfF+ejytLrAwMUw72yOrtsafqB2YD7/P6
hAoE143PnsP7mt2kWONPLDooAGwSn8emtAPj5dNTeh9ONiycY+jJZKtXusP5bAGP21NzN4nQ
8ccrYAgYYX0MUSnoXU73GMD0C/VFXexCOrloc6fH+7Zg+iTNN5ntIMU+xJrCMqCd+qUwCHWK
+WaSgqQzUE+zqKpTmpZ02i1crZ2gDB3XZSRKUSsNKP8TlgVbGvnCr7Qh/HgYYeGdfznLIrCC
/Zw+Yr7bWRM699OrewrTVwONjyVvZ7GccnLJeO62iUVs1nPDRn+GfYjSteGsPpAl8a+mCxKF
6bxd2wbR/BxVaseoVuJjbxc9Q8D+onyJe9x3KlLegMs9ukMHddrNejFtLLNAgzJVj/hi4OHv
D6zLk+EBVXPJy0uUoqlzevJLmiiuBY9kYLqHbTyAqv0uxIR4yDu+kq581uRxHeKPt+S73eCA
zpwf3CE167EFeDoa+Mu0kghkEji8zZ0HbwYjd+ZW48IqH/lE3cROJ2lIhqcWnBy2n+saHAWG
nnkZsDl6ZutI4JP83G2gdG1l3cF7J8TvI9NIJFFgTo9PNiKTO3NdglZFTlTMFWPoKrI+5Vg7
MpaPWYpaKKqCgTtXsN+MExQyJl/JDGjDTxSDpdd+SDi1BjrEyVlNSmeQg3J5epyPvBdQyMFo
M0qT0lpeBLYNZLJ+Vbv91mNeNmcFgjS37JPgmeWagzrBZ6pvkLHzowgxUG9yoFKn03qXryxH
3b9BHAqGKxcyJ0WG4nKAND4IJwm6Jo2mHGeiL9z2iJ+mA60/3Qb+wd3Ct1hEGSDxijuCSPf/
fTJwNPrrsHpdWSnv3LmKut38RMZUxqQZoM+tPymlD8in96XsD/rnjW/rZcX8coDObxzVVtnQ
P+289fFOuuprKfmA7eLZEqg7rcKvJ/y6WYUo0bB7p1IcI5T8wF6iLOr/gjMi5lPIYrHv/0Ul
MwXlNyja1/bXVhMuUpmcTkv+iCNIwgh2AFEzqS/uoUmYyy+6cOLBXKDrnZ4M9BCMeAe92SXi
25PR0kuqd1K5wdyWDWPpQXy/nrT0fNB+6an40E0fv/sLHC6NF9MxwqawHRwSOTW0TG4grPro
F92/672JspkHNGIcbcxt1I8zn5bjH6qYLe7Q0E/A71yYERBE1bjE6JXWgq8aob4eexadI637
dNUxzj8FY0Wo8DzKzymGzXHFvEYaEzWU+hVB3atxITC9RK2halF6Y49uMlnXQedoqP6KoskQ
Nvl+M1orzjMaL6VRjLng7sG5/ZKLvt+jc5WD6RUbhczN4bcZCNMzyutadHAEF4r9OKvppJZ3
W7W/voRaisDCfXEEAJpB1z94kSRPhCUapP0CkUKoppol3pT1D7Sw+FDo0UI3ygWvk1eMSlAw
oF7wQliV8uNzDQZXCag733PiWVhvTEo8ReSbgVMDWEN9LvFZaEDBkadt7+EwALaFbqaIpQcd
Ebni2AbNcJeHORi5/+GVgDhZzWU5EROstAOjsW0xLHikAcOQO5Xv01JBJNqwLcHbMkX8MiRG
S9BZG1fW22OEz2g0OMaUVPZ1pXgFkaAn/Ayddoci3ChFP5Uqwlk42NpZQNAQI+1jlQnFPQx6
HHddocEDjgWo+1QEjXN2oR+JsVLOcn6Q333T9ct0BzuiJufrSSjhWV4F6vAYFMKgu1uTqdQl
iW/TF/B3HjVB5HTMJns9OjjuJwxF0+LBQV2V4qmAm8VIoDHJSNiJdbXz59vdHmcasS4HkYrC
Cmno+etbz99YBnGZEOBUbvzDf1z4ZqBgfM4NUAlW5hZ0oMor6j9MlZbJWoT/hAsDJy6vlAfK
pQDMXDjE8QzdU122lxuwTeATzOfo2kXwraswhpCY7gdJQhM97L/Tdi93g4frfXYECRx0kUWB
c5rsLKrIpaJisybA5fOpfNCN+MxA/IeLqWYQpfTZpF7mEWnWKCQWsuj2swWQmBx1Eb9WIQMS
QrawsEeIbWmn5dtmTMYgkF5Q+kpTY5QH9r2d5+74AxPONQuF70D6IYcQRy3yvPhYOvyzfRvL
ZOYhGWUQTbbrX8q9A7XtT3a0Ypi2Srrs5bPm9oykriTfHz9vp/05obkTYiJa7xnJh3m/Hx22
nxUSmPDKspkJBy6PBrGixBQGjO3K8lM7+fGUfgdMhtoi6rgXLxrlxEtSlXbySy0CgUsVuCJz
qYH0ekhZXuo+rVcan5B5GNHeE880M2a+nYTBNBFmVMKLJurKie0BVxfT1L1WBkywFle6Yfjt
SjFPhQkhThouUa587U7nsZNrZftPYmWFJWGL9QUY5qrcl9jIqMsmlyYZnhZxbkSo5uzvkaTw
rox2XohLfUOt+QlLRaFsdtWLhUsReAX7jfnXJm++mx4IxPEfksXjJn74TQ0ga4cVuZ9iC1H+
6lrW/BTBdYYgdj0iu7JO0LxUG3o1mkFCEShnkb2wmVeOrYJVKhBi2/a/4wHOVeuPOs3qFFEw
YTyVm+w31W6AgaOx86yThuQmdPrqAsxaOfnmxx2a8BHro1ghejc2d3p6G51Qu1/18vdkkrXe
UP7+1uXXQcvdEQc0uarWn1D9o7LlF6gw/aRUGCcJSiT1pYMJgKJGn/TSjsOSxTW/hLjRDFeW
w01Q2RrtQNCvqTyyaxvK8O8DQiUe4iTUCo/VKl3EuKB2lLJyRYZYMDl5FJJplcn/Ous6MTpy
F2rPpJpKatTa/E6tCnyCvhG9/knplSH7iKRzcUHKV/JkxQhxj+HSw16x9CXOCPcXjYKYkVOH
LChbJ7WTtJLWtGM2Pw6P6J3keztnyXC4gtLEPI7zsLS05Twgj8vkowG3lPQKuXJDqeagnZGx
KWZVJHimRooM+qAtQ3UnayMYrDdJGUpdp3q1KwUfy4iyw07jMZn5AG7+8etqpLXai18/M2is
eJzP/Yhax1HwmnBVdbh/g4UGZJHuElu0aOStczcSx2sAESaTxGj54RsvMfORl0KQ1Ut25nM2
ipWvj3/mttCzVT+KUIOlI3/CXk6pEAVfYh9bSbETl0DBSuEXZerPQN1uTjHPv0oeRLayWiz4
p3rM0nM/W9yu7dBOzdcBjaH3jwUmSFaUYRuXVNJ+GIbzzeJdYFkZ9JqEUGVvhd53TiSWWmBS
vwxEYmUfQIKpvP5261j/N+ImElc2ZmJaLbBQWOSAZ2iZAuVwxiGftW6xPWqv6j8GrHjmGcMG
7yLlYEEHyMssYM696bAUZfJeGD3tUNZts6Naii39/uvQFF4N+3kk885gfTHaa74pZIt5QNvE
vGFHmbi8QjoG84k0YyafU9Op7gvZGj18q3fzBxtDsZkSKNca9bXsjX8CXnO3PLI6uMMOH8nu
shBun7OamEYcxocZcZBen5r2v9DDkQ6mVEMvC3Lq6rhqBrCYYLHm/lUvKMX7pjhB6B4r72b4
FBqCXGiir0z0AHfElDnbRpIPBPFmtMl+ii/vmd2jPvSdygAKsDyxuYd+wihK+EGKT6QU9ysA
su9TJFGsZGevblPUqZo+Pxc1QcDk1BxU7XBHKHc2TF5G624L/i0KfHfHYc6CayH5ABP/2bdb
TTMvXY3AKlZBNxR7M6dfA/qvDx8xqTsdrggXTP6jZlRKpPNuckbWK8B4N1TBZ5EdTXYvKX7J
DeAJGpaMy8+/1q8EbQvRPPL8xwXOzfEGhD506H5tlKjr60gBrZcDizm69wvMlcuh64TUxq4k
zVTVU4Khz4nTkF39vptUUUkI8pzGlliGKDSQYsdvTypxGUVVCzyOHriYPgoYODwG9VJ5H/7e
5ycNvNslFJ8+X+Fjd+OWOM4MKnv9jsjHlBDvjsRDf0VAfCGaNl3aTu2lChRPtvG3nIQtMgSy
WGp+l4ZNMspcqFY/AOKLK6zQT/Jl9I3O0y1n+ogITo15wZGRSOfjcBzW+6PINGF/ibdBh4nK
a6CfVmgTweTtDUBp16gz+P2I9GL2I1syT8Rr5sAwf7PdEa7uHVFUtMBDHbIrxXnaGQdl+rBx
ARAUOf0OzV3Z8V2n4IN6zwuo+rqdUbiI6Ygrr8unCWFCHJbeI4pnunnIhX+NBwlb+W0PHtWJ
zvGKE4CDqGauvxTyvL9Vm3fMpHpTKSlpdMpF3afxrE8a4x4akIQ+4mHR8Uahr2mS1z21Q6WR
+4/POgvCdods+RyIuB2qXnm2BBDZm+cVy84BRSVIA/KM+oxCYs5YFffvCr4pxCHPNjnfocJU
UON99+AoUOzUU6146kP585fsf9WAdq/Dp0WkXzcUXZcyoKC6ulpv8yhjlU4J9MbuSO0hJ+O7
RkQyhU9UVnKdUb1mZYTQfFPMjphN3O9EZLQZuGb42ZkKbm1NfZt9ZSjmxvjmTlQR+43a25Km
GqS8LgCxM/+k5gtFYRJcVSvRgAdN7TVnngx3NifsSm5MFHogrpgAa1km77XPhUu+YPyBRNYu
CYJIukzAnGCZLziq3/+tuzMMc7Fcr0oRSuph2FMeIo0ot6vQBTf2+PWLsjK6FyrSPx+1ZKJo
C4L51piZTacRf0ymG6t0UHym/5PRyca2wAM6aOlgLlmh582otkKzPwnj2Bt1rtlCNHQhSl5k
3aF7E7wTNjNzK/JqWub6PaHPSoQcP+VSZeWhe+yXyTm/ktqg2MIqKNxNRmgKikB+gmYM8WoK
TTKRZZ5RI3t+SuH86B28icuEB/N41YEUF9j1MKM+PIiW/Pdq4wc/blSRk4GuQVnrhKvcZrxf
2U8PQDE8W47ZmakIoSrUmTJe/Q3esOKPqdBE3jePRxkJJDKHI7PgVt0NpN2+m5/63kEk42Pr
W5eCWLY8Qwl4dnb+kaB1xLl4gouiVjw4FpmY5Y4FQhJdq3tKhLjN6BHCE9O99q7RdLpfbjBR
EciZQjDrmFWiHENEOVpMDsQQmNH3vdUh5xwzbvg3U2hNmvrVJUdSDYHuT5rAKGIfHIt+swJy
mt2VARwyOhrdKEXzKw4VvztB+lPRSTW5HHsFvKH22RFA+Q66FCC9MYKALgs8aqZKb2OmEAr2
LKxQs6v/WDvWytOOA5R2wtbWNsKmF86tEzw5+ro7tz3+CuYo7L+ZGqaNcbcJKwflB3WFClrL
l9LJbil6RVzs/hl3e4TTIiVJqL5OQ899F47NY9/0z9FOb8UHXZaNf7wPtN4C5FKSmUjigZnq
qSidpyGFuAV61zjezJI4JYsu+//J8mHeIwUotsN454Ycmd0Yr68I2ySOIkC04Gvf7sN7Q1n7
pDdavtz5Xqfriu3d6L57JFOeO90PZ5b+cGjzetTwc/wgZZDBRyZH8HFTFCwTZDfsktnV1Mj0
6swcscG/HpxOYzUISWIowknMSKLO+EMfO2iemnE+RmxNqptOrqzuA8p0vEoky19nRdmwVpPe
CNzFlFtmroIRYiAoZEJ7Ez0wC1ZGgTbWNZTGK8rpJqGlHhEJHl5iGP5I3WpcHsXVIrGZqaAs
PYfqA5mbZr7xxwtqUqiWN5kqI/w4jvFpRII+R9qLFqXJoJiFgnAhEQpaTqjMwhD4hFRh5Ne8
URP+5r6fNkTECylUGqkR1mxuZOflbojTtjHJbOH9DWeBGCBuTxxroydx0RKI3CWEXikAMgS7
MMjFG0Varqlxx4i0OHEoyvUi3YO9FxoY8phWEk3lPD2j9/ki/noNUQccty7CROAv8WzcNRfV
lPHMtg8bz/d80c0WYClU0WAQ42sjaMtzvxeDKbrQRROrEJTqfiVlwrLI3dvaVolJaTp8NNPB
sfEaMeC+3BlB7DF6tH4WpXB5ZmjF9HuQAmA37aD0SMRcyDnS3CVjgjcwMH/BodBB9aD+MNjx
pQjhJKX7xss2+R6v1DgCW1QvoCgZNZzG8RkjgQaFRVE0qVl7bR0tVxYSh+VVigYxVLxdrISH
0trcApPzVgL2Cj5hIitVypsf+cUJcvozxl0/grY0k1yZzBvRMdfxYM2skN7DBfSR1mR/lY3q
V4i5Qo4xbFSsQYh29Rxokx4J244ATaHFgaEmNUgoeVEJXog89VHbzeYQy0PFsmENDVkJutxw
VxxSZcwG/h7JG61iPWBbSX27I6a2EjC2onMkO3YyvZQCOFGtGOJZqg3zEV+tiiV/6vNgn5hF
Dm6ov19SZjnA284JKJZT8Y9PbZ+Ul3QvEq2UMPhAKwPxmb3/9D1L3C7Qa5dPeQMDYsSAJbjd
U/jMzH0i7wun34aiarXjtb257zxRHzFFSYGJ4viUlXsgyRfsCsUojCX1n20t+geXkOh30AkE
xG4rGEV1zwh0ar1AJehbSi09un62kF3Jd9g4v/KWiJ+RZ3C61RGtac7+pl7ARe7sBLVYeNYG
hHJgxjgBje5KGs1qEsJoE7f+DpPCN9t9W7mikG9qUTALHf1soNW3pMnuvM41s8p5TgKMpMsU
O6CTXkH7E7TJR4xTddTVnS4MzhVEhynllRj5F5/qxSzEZGcFVLNJlalutupVGkCe4+q6pkl4
xpLeO81E8jE1syCUc/8pfyIqtceyyyIBzSfZcjNPcfCQrDfe4DN2AncXTq76SphrJKZH4Ha4
NBUaNgY8+g1/aUMAPtgV4moJYNwqYuZBI01EnvdyhEfd7WiapcHisLg0BfCcp3jrae1c7TpP
+6KL8T2w/x7T5pfu6TJlbitZ2p0frRBwctfIgK4PnkKZ4giP8BnhXaFtY4ZAt7pofDjiSDnn
tNCqdwrK5g+ignXeUMLYbvP1/vFKbsk5SOaSMiKhIABVK4MVBmj62xpGG0mpHgdiycg8SjqY
EaXW+skQ3XTx3zOMsOiuLYxidxFqY7QgKHkHZoJS+PrxloXDYZcRvxXWmjest16/Zlt5mwFz
hbENDnXTQsEUQHc0P3AZPTfqxDPv3Qg8jW2Q+rVeJmalwFgiXYj+f/W7bB3guH68ThdBatE+
ZR1/0TkzB6izi2VE2iWW7HnG8pcZ6bDtujeVATf8L91wvM7gqyvgJOGbyEUdTQPz/LH54Lqx
92BSFi2xaRhZGCIqPqE1svxSq02QNotY9GV2oTYaI+1METkVkHApUmmQpTMHxAwQJO7wD3rI
WusVGsQNBA2f+6sxNcs7YzBUeX06oGrvQd9MjsKbr2GFLoiz+sUN3iEcj65JIXgp9BF43gOH
2epSFkEGD179LQV8yuAs84pkm9AbWpe5gtGJyARNhAccdhA/22E9RspnhTnrE3j9RkmPDEiH
5FSC2bt3sD1ZaW6WgYyfajnMOABWSB7Tk+2kR/Jx07fo+1/HLna7DSPL1AiMPTba6BIH+MeC
JDonwjzULQHU1jnWHrlPBRIpF486nvSbix9ZNzZ5TZ3dIi5kIxFZUfJS6PE2iTPwDwYAi5/R
fQ+NMp4kCGLX5OYm5pMx6z0+U7tWl0og31pOzntnRU9Qu05CEEocq+z6Pwp9jNR62/jNGMg+
z8YmS8TER5TYSllUxdQTlb1eQ3ApBinonSEMnU2SicbVwV43hIdpUZjbqP9sHCIw5mlxwv7E
QxZWnTIX8bRF6gQSBf/24SR5jKIPmyiLLyDmd3uy5IjlveAlBC7PsMOekXIAdFOeiV+U/ws2
WADsR/h+WMqcV9euxzVASrA+uObMjFKTElNdeyltrbQ+h6NbP70p1FGCNT6aBn9YqgXQgBaf
aEtZI1EskKF7qIg3OoKxCx4VXiwSyRKZpWqV3BwxLHe0YReHScEwKugfjp7rxoHi6RE5gMij
sU7fv8eaF/b3mf6DnMMb/PD4FD7PzBnUROPq4LxQw0v6sKu1swN1Ll84gUXfEEBUOVo9jlcp
Rkjmo+ozMwYUrsJZ7tWOTVrI7oTiWuKaK+nAaMciD6nesXvMtmfGS3W68BS4Oaa6/kMcYsTs
APjv/2NqlbQLOY+5MluUe+x6rogsvB5g48GjesLcq8rBZGXCJz36M7WpWnHtKk6PV7Mm3ryu
y/3923JhS7uVtzzYgbfi78kIc8CL9X8g6VLvniGU+Q7Zpd8cbnkKgCX5LBXdIEl9GX6rDE5K
bZ9Smk3glpoaAPbNNYwxfWF44ntxTpwPR5W0lVrKS4i5V/8ZuN6BbAdCIgSffGwD3aWCC+Vi
I+r/k/BnFegMQOELWArPjgnbzXSrlgNoOl/7hSfG13xoi+pbv5M9C0Nt+YjHp3JV6qrvN3CT
+5WS6V4lbLMboX/lIHBedGF9Wq9zBd0zlN66hKARaOSkgSnW1KhsdBFRvmzDgkyyCg1wMS7P
zRebS9sB2zTKJlCdT/iWxBcBguSDru9+EXPIpbgyWWDqf9r2FQ8prTmkb2TqvPB77YpSS9Dq
iTdYLu2gCTs35y2Mpt5rJx3uB0NsLM/uCX3u+VnbdCHpZlJiFronzed3g3UUXvx3KUyeGM7J
Z+Pn2v3gx/lOtjZTdtJ1K6pG/Pa3bhQZ94Jwt95l6BF5giIzLyQQ2nQqtv48FFJEdT6Y63h3
nX+t07X3UICcJUMHBaJvGp4IItnoKGfkAmm1SrUNyO5yySaUojdK/9bOqzggRqk8sBpuNUuO
5ZuWkyUIw/ZgnGgWauvyrrxWicKU83rXb6cwAAklnScoTqWGoHJtz4Nwc5vlhsjZP2d+YONZ
5607BdweF5YkLfnKBBHacI5Aj3jiBt8Fv9x4cvFKFH0+aGDMmEHJ9IDo/u9Q1+Q2w0FRrDer
Zbu4yccu2Kl9Uez4MdIJ+9ydeiKvKZeUvJfpclYfasvf1nnuWCxMsw0JtGkKT1+B/iAZYeek
eKwIBZ5QvjDiT3MqJZSYVeHiw5skwXnebWUir7rfesyoot7Fq7Guw6iImBXg0QW7D5s0OBnU
JsWl4zhMXEOsgL2/Cd3hQb9BHLwMsjW4NirImLJ1zYKPWAgE1zr+BGOzBRA89as81kDDSu7S
8EpSnY4GSjCXEBImWl+doEO1VRnGKORFrfUjWK/v8xhDrjY3Q7Vi5QqXVdsuXrHkOAgRqQPH
yY/dKtETtlxYU5cwVoOnsEuaAtF/wmBE+C1/F4hlEyPT53Yk2nkX4mNdAOZYNcawtrADpIZx
05pzFI/BMfByfAUV1tf9pt4Jnnk0mVP60H6mQVyGyExLKqGM+kA9agicw4str/q/ajXGaa4Y
FZ40gVp79ib5ri59rTm5rkYu1O8zU0fCan2s+51arpuG+qV+YdM5l0yFc5dKjAI11EfZGdwM
GLCmW+LXrCyoRsmaV8vxa/0EHwrcshNRpVHITkF85htPR7Y7zjBHHRQc6ojNKGCDf7fsvtq1
eWgoOWealb+sjKy1aNYQmLv3S1Ee1BKxTxIBs0yp3/HraGQHuUNpqcZjnsZKQrvOml7WNsLT
Xhi8e2EcxsewiGr3o9UpRBUIxOFVK5n6EoWpk7XKobFs3Q2GNasLPJkW+Z4ZkComKTnCJ9Rz
JJ2rh4j+BcLL9C/CAQr0YpmiXpkjcvkg3/rdD1KLugmlyFVdHtVYCnguQrdQohvE3nqDKFXF
5+oQs/JZX2D9POpahwv7dN9W/hfrp2EHcAFWABkXSUXsh36hIJ6/6VSC1Dh+X/DyJAak7g35
USiqycLDSkhEyp5w3WwbVVQcaIv8QhBFY2Uau/Q0QCY9EfJhV8HnIeeABy/MWvnqrTI4a7Sn
qfXehF7L4i/IMGPA+PC/dNtkkG8v2U+2+g0P4kKGRQodBf2DXsso63HeVL2r/w7uShPqnT3L
BDYP82L3PPfowzTmQCmPtNGQqeTHng==
`pragma protect end_protected
endmodule
